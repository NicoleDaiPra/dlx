library ieee;
use ieee.std_logic_1164.all;





-- ADD BITS TO ENABLE THE SAMPLING OF RS AND RT IN THE ID/EXE STAGE REGISTERS
-- BECAUSE OTHERWISE THE STALL UNIT USES THE WRONG REGISTERS (THE ONES OF ID) TO DETECT FORWARDING







package control_words is
	subtype cw_t is std_logic_vector(61 downto 0);
								   --  ID	       ID/EXE      EXE               E/M    MEM     M/W WB
	constant rtype_cw 		: cw_t := "00000000000000000000010000000000000000110001101000000000001000"; -- because the signals are determined using the func field
	constant bgez_bltz_cw 	: cw_t := "10000011110100000011001100000000001000110100000000000000000000";
	constant j_cw 			: cw_t := "01000010110000000011000000000000001110110100000000000000000000";
	constant jal_cw 		: cw_t := "01001110010100000111000000000000001110110101101000000001011100";
	constant beq_cw 		: cw_t := "10000011110100000011010100000000001100110100000000000000000000";
	constant bne_cw 		: cw_t := "10000011110100000011010100000000001101110100000000000000000000";
	constant blez_cw 		: cw_t := "10000011110100000011001100000000001000110100000000000000000000";
	constant bgtz_cw 		: cw_t := "10000011110100000011001100000000001011110100000000000000000000";
	constant addi_cw 		: cw_t := "10000011100100000100001000000000001111110001101000000001011100";
	constant addui_cw 		: cw_t := "10000001100100000100001000000000000111110001101000000001011100";
	constant subi_cw 		: cw_t := "10000011100100000100001100000000001111110001101000000001011100";
	constant subui_cw 		: cw_t := "10000001100100000100001100000000000111110001101000000001011100";
	constant andi_cw 		: cw_t := "10000001100100000100001000001000110111110001101000000001011100";
	constant ori_cw 		: cw_t := "10000001100100000100001000001110110111110001101000000001011100";
	constant xori_cw 		: cw_t := "10000001100100000100001000000110110111110001101000000001011100";
	constant beqz_cw 		: cw_t := "10000011110100000011001100000000001100110100000000000000000000";
	constant bnez_cw 		: cw_t := "10000011110100000011001100000000001101110100000000000000000000";
	constant slli_cw 		: cw_t := "10000001100001000100001000110000100111110001101000000001011100";
	constant srli_cw 		: cw_t := "10000001100001000100001000100000100111110001101000000001011100";
	constant srai_cw 		: cw_t := "10000001100001000100001001000000100111110001101000000001011100";
	constant seqi_cw 		: cw_t := "10000011100100000100001100000000001100100001101000000001011100";
	constant snei_cw 		: cw_t := "10000011100100000100001100000000001101101001101000000001011100";
	constant slti_cw 		: cw_t := "10000011100100000100001100000000001001001001101000000001011100";
	constant sgti_cw 		: cw_t := "10000011100100000100001100000000001011011001101000000001011100";
	constant slei_cw 		: cw_t := "10000011100100000100001100000000001000000001101000000001011100";
	constant sgei_cw 		: cw_t := "10000011100100000100001100000000001010010001101000000001011100";
	constant lb_cw			: cw_t := "10000011100100000100001000000000001111110001101100011000111110";
	constant lh_cw	 		: cw_t := "10000011100100000100001000000000001111110001101100010100111110";
	constant lw_cw	 		: cw_t := "10000011100100000100001000000000001111110001101100010000111110";
	constant lbu_cw 		: cw_t := "10000011100100000100001000000000001111110001101100001000111110";
	constant lhu_cw 		: cw_t := "10000011100100000100001000000000001111110001101100000100111110";
	constant sb_cw 			: cw_t := "10000011100100000000110000000000001111110001110011100010000000";
	constant sh_cw 			: cw_t := "10000011100100000000110000000000001111110001110011000010000000";
	constant sw_cw	 		: cw_t := "10000011100100000000110000000000001111110001110010100010000000";
	constant sltui_cw 		: cw_t := "10000011100100000100001100000000000001001001101000000001011100";
	constant sgtui_cw 		: cw_t := "10000011100100000100001100000000000011011001101000000001011100";
	constant sleui_cw 		: cw_t := "10000011100100000100001100000000000000000001101000000001011100";
	constant sgeui_cw 		: cw_t := "10000011100100000100001100000000000010010001101000000001011100";
end package control_words;