library ieee;
use ieee.std_logic_1164.all;

package control_words is
	subtype cw_t is std_logic_vector(52 downto 0);
								   --  ID		  ID/EXE     EXE                E/M  MEM    M/W WB
	constant rtype_cw 		: cw_t := "0000000000 0000000000 000000000000000110 1100 000000 000 00"; -- because the signals are determined using the func field
	constant bgez_bltz_cw 	: cw_t := "1000001111 1000000110 100000000001000110 0000 000000 000 00";
	constant j_cw 			: cw_t := "0100001011 0000000110 000000000001110110 0000 000000 000 00";
	constant jal_cw 		: cw_t := "0100111001 1000001110 000000000001110110 1100 000000 101 10";
	constant beq_cw 		: cw_t := "1000001111 1000000110 100000000001100110 0000 000000 000 00";
	constant bne_cw 		: cw_t := "1000001111 1000000110 100000000001101110 0000 000000 000 00";
	constant blez_cw 		: cw_t := "1000001111 1000000110 100000000001000110 0000 000000 000 00";
	constant bgtz_cw 		: cw_t := "1000001111 1000000110 100000000001011110 0000 000000 000 00";
	constant addi_cw 		: cw_t := "1000001110 1000001000 000000000001000110 1100 000000 101 10";
	constant addui_cw 		: cw_t := "1000000110 1000001000 000000000000000110 1100 000000 101 10";
	constant subi_cw 		: cw_t := "1000001110 1000001000 100000000001000110 1100 000000 101 10";
	constant subui_cw 		: cw_t := "1000000110 1000001000 100000000000000110 1100 000000 101 10";
	constant andi_cw 		: cw_t := "1000000110 1000001000 000001000110000110 1100 000000 101 10";
	constant ori_cw 		: cw_t := "1000000110 1000001000 000001110110000110 1100 000000 101 10";
	constant xori_cw 		: cw_t := "1000000110 1000001000 000000110110000110 1100 000000 101 10";
	constant beqz_cw 		: cw_t := "1000001111 1000000110 100000000001100110 0000 000000 000 00";
	constant bnez_cw 		: cw_t := "1000001111 1000000110 100000000001101110 0000 000000 000 00";
	constant slli_cw 		: cw_t := "1000000110 0010001000 000110000100000110 1100 000000 101 10";
	constant srli_cw 		: cw_t := "1000000110 0010001000 000100000100000110 1100 000000 101 10";
	constant srai_cw 		: cw_t := "1000000110 0010001000 001000000100000110 1100 000000 101 10";
	constant seqi_cw 		: cw_t := "1000001110 1000001000 100000000001000100 1100 000000 101 10";
	constant snei_cw 		: cw_t := "1000001110 1000001000 100000000001000101 1100 000000 101 10";
	constant slti_cw 		: cw_t := "1000001110 1000001000 100000000001000001 1100 000000 101 10";
	constant sgti_cw 		: cw_t := "1000001110 1000001000 100000000001000011 1100 000000 101 10";
	constant slei_cw 		: cw_t := "1000001110 1000001000 100000000001000000 1100 000000 101 10";
	constant sgei_cw 		: cw_t := "1000001110 1000001000 100000000001000010 1100 000000 101 10";
	constant lb_cw			: cw_t := "1000001110 1000001000 000000000001000110 1100 000110 011 10";
	constant lh_cw	 		: cw_t := "1000001110 1000001000 000000000001000110 1100 000101 011 10";
	constant lw_cw	 		: cw_t := "1000001110 1000001000 000000000001000110 1100 000100 011 10";
	constant lbu_cw 		: cw_t := "1000001110 1000001000 000000000001000110 1100 000010 011 10";
	constant lhu_cw 		: cw_t := "1000001110 1000001000 000000000001000110 1100 000001 011 10";
	constant sb_cw 			: cw_t := "1000001110 1000000001 000000000001000110 1101 111000 000 00";
	constant sh_cw 			: cw_t := "1000001110 1000000001 000000000001000110 1101 110000 000 00";
	constant sw_cw	 		: cw_t := "1000001110 1000000001 000000000001000110 1101 101000 000 00";
	constant sltui_cw 		: cw_t := "1000001010 1000001000 100000000000000001 1100 000000 101 10";
	constant sgtui_cw 		: cw_t := "1000001010 1000001000 100000000000000011 1100 000000 101 10";
	constant sleui_cw 		: cw_t := "1000001010 1000001000 100000000000000000 1100 000000 101 10";
	constant sgeui_cw 		: cw_t := "1000001010 1000001000 100000000000000010 1100 000000 101 10";
end package control_words;