library ieee;
use ieee.std_logic_1164.all;

package func_words is
	subtype fw_t is std_logic_vector(62 downto 0);
							   --  ID	       ID/EXE      EXE               E/M    MEM     M/W WB
	constant nop_fw 	: fw_t	:= "000000011100010001000000001100001001111100011001000000001011100";
	constant sll_fw 	: fw_t 	:= "000000011100010001000100001100001001111100011001000000001011100";
	constant srl_fw 	: fw_t 	:= "000000011100010001000100001000001001111100011001000000001011100";
	constant sra_fw 	: fw_t 	:= "000000011100010001000100010000001001111100011001000000001011100";
	constant jr_fw 		: fw_t 	:= "010011011101000000000010000000000001101100100000000000000000000";
	constant jalr_fw	: fw_t 	:= "010011011111000001001010000000000001101100111011000000011011100";
	constant mult_fw 	: fw_t 	:= "000000011100100010000100000000000101111100010000000000001000001";
	constant mfhi_fw 	: fw_t 	:= "001000011101000001000000000000000001111100011001000000001011100";
	constant mflo_fw 	: fw_t 	:= "000100011101000001000000000000000001111100011001000000001011100";
	constant add_fw 	: fw_t 	:= "000000011101000001000100000000000011111100011001000000001011100";
	constant addu_fw 	: fw_t 	:= "000000011101000001000100000000000001111100011001000000001011100";
	constant sub_fw 	: fw_t 	:= "000000011101000001000101000000000011111100011001000000001011100";
	constant subu_fw 	: fw_t 	:= "000000011101000001000101000000000001111100011001000000001011100";
	constant and_fw 	: fw_t 	:= "000000011101000001000100000010001101111100011001000000001011100";
	constant or_fw	 	: fw_t 	:= "000000011101000001000100000011101101111100011001000000001011100";
	constant xor_fw 	: fw_t 	:= "000000011101000001000100000001101101111100011001000000001011100";
	constant seq_fw 	: fw_t 	:= "000000011101000001000101000000000011001000011001000000001011100";
	constant sne_fw 	: fw_t 	:= "000000011101000001000101000000000011011010011001000000001011100";
	constant slt_fw 	: fw_t 	:= "000000011101000001000101000000000010010010011001000000001011100";
	constant sgt_fw 	: fw_t 	:= "000000011101000001000101000000000010110110011001000000001011100";
	constant sle_fw 	: fw_t 	:= "000000011101000001000101000000000010000000011001000000001011100";
	constant sge_fw 	: fw_t 	:= "000000011101000001000101000000000010100100011001000000001011100";
	constant sltu_fw 	: fw_t 	:= "000000011101000001000101000000000000010010011001000000001011100";
	constant sgtu_fw 	: fw_t 	:= "000000011101000001000101000000000000110110011001000000001011100";
	constant sleu_fw 	: fw_t 	:= "000000011101000001000101000000000000000000011001000000001011100";
	constant sgeu_fw 	: fw_t 	:= "000000011101000001000101000000000000100100011001000000001011100";
end package func_words;