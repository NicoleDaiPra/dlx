library ieee;
use ieee.std_logic_1164.all;

package control_words is
	subtype cw_t is std_logic_vector(57 downto 0);
								   --  ID		   ID/EXE     EXE                  E/M  MEM     M/W WB
	constant rtype_cw 		: cw_t := "00000000000 0000000000 00000000000000011000 1100 0000000 000 000"; -- because the signals are determined using the func field
	constant bgez_bltz_cw 	: cw_t := "10000011110 1000000110 10000000000100011010 0000 0000000 000 000";
	constant j_cw 			: cw_t := "01000010110 0000000110 00000000000111011010 0000 0000000 000 000";
	constant jal_cw 		: cw_t := "01001110010 1000001110 00000000000111011010 1100 0000000 101 100";
	constant beq_cw 		: cw_t := "10000011110 1000000110 10000000000110011010 0000 0000000 000 000";
	constant bne_cw 		: cw_t := "10000011110 1000000110 10000000000110111010 0000 0000000 000 000";
	constant blez_cw 		: cw_t := "10000011110 1000000110 10000000000100011010 0000 0000000 000 000";
	constant bgtz_cw 		: cw_t := "10000011110 1000000110 10000000000101111010 0000 0000000 000 000";
	constant addi_cw 		: cw_t := "10000011100 1000001000 00000000000111111000 1100 0000000 101 100";
	constant addui_cw 		: cw_t := "10000001100 1000001000 00000000000011111000 1100 0000000 101 100";
	constant subi_cw 		: cw_t := "10000011100 1000001000 10000000000111111000 1100 0000000 101 100";
	constant subui_cw 		: cw_t := "10000001100 1000001000 10000000000011111000 1100 0000000 101 100";
	constant andi_cw 		: cw_t := "10000001100 1000001000 00000100011011111000 1100 0000000 101 100";
	constant ori_cw 		: cw_t := "10000001100 1000001000 00000111011011111000 1100 0000000 101 100";
	constant xori_cw 		: cw_t := "10000001100 1000001000 00000011011011111000 1100 0000000 101 100";
	constant beqz_cw 		: cw_t := "10000011110 1000000110 10000000000110011010 0000 0000000 000 000";
	constant bnez_cw 		: cw_t := "10000011110 1000000110 10000000000110111010 0000 0000000 000 000";
	constant slli_cw 		: cw_t := "10000001100 0010001000 00011000010011111000 1100 0000000 101 100";
	constant srli_cw 		: cw_t := "10000001100 0010001000 00010000010011111000 1100 0000000 101 100";
	constant srai_cw 		: cw_t := "10000001100 0010001000 00100000010011111000 1100 0000000 101 100";
	constant seqi_cw 		: cw_t := "10000011100 1000001000 10000000000111110000 1100 0000000 101 100";
	constant snei_cw 		: cw_t := "10000011100 1000001000 10000000000111110100 1100 0000000 101 100";
	constant slti_cw 		: cw_t := "10000011100 1000001000 10000000000111100100 1100 0000000 101 100";
	constant sgti_cw 		: cw_t := "10000011100 1000001000 10000000000111101100 1100 0000000 101 100";
	constant slei_cw 		: cw_t := "10000011100 1000001000 10000000000111100000 1100 0000000 101 100";
	constant sgei_cw 		: cw_t := "10000011100 1000001000 10000000000111101000 1100 0000000 101 100";
	constant lb_cw			: cw_t := "10000011100 1000001000 00000000000111111000 1100 0001100 011 110";
	constant lh_cw	 		: cw_t := "10000011100 1000001000 00000000000111111000 1100 0001010 011 110";
	constant lw_cw	 		: cw_t := "10000011100 1000001000 00000000000111111000 1100 0001000 011 110";
	constant lbu_cw 		: cw_t := "10000011100 1000001000 00000000000111111000 1100 0000100 011 110";
	constant lhu_cw 		: cw_t := "10000011100 1000001000 00000000000111111000 1100 0000010 011 110";
	constant sb_cw 			: cw_t := "10000011100 1000000001 00000000000111111000 1101 1110001 000 000";
	constant sh_cw 			: cw_t := "10000011100 1000000001 00000000000111111000 1101 1100001 000 000";
	constant sw_cw	 		: cw_t := "10000011100 1000000001 00000000000111111000 1101 1010001 000 000";
	constant sltui_cw 		: cw_t := "10000011100 1000001000 10000000000011100100 1100 0000000 101 100";
	constant sgtui_cw 		: cw_t := "10000011100 1000001000 10000000000011101100 1100 0000000 101 100";
	constant sleui_cw 		: cw_t := "10000011100 1000001000 10000000000011100000 1100 0000000 101 100";
	constant sgeui_cw 		: cw_t := "10000011100 1000001000 10000000000011101000 1100 0000000 101 100";
end package control_words;