library ieee;
use ieee.std_logic_1164.all;

package control_words is
	subtype cw_t is std_logic_vector(54 downto 0);
								   --  ID		   ID/EXE     EXE                E/M  MEM     M/W WB
	constant rtype_cw 		: cw_t := "00000000000 0000000000 000000000000000110 1100 0000000 000 000"; -- because the signals are determined using the func field
	constant bgez_bltz_cw 	: cw_t := "10000011110 1000000110 100000000001000110 0000 0000000 000 000";
	constant j_cw 			: cw_t := "01000010110 0000000110 000000000001110110 0000 0000000 000 000";
	constant jal_cw 		: cw_t := "01001110010 1000001110 000000000001110110 1100 0000000 101 100";
	constant beq_cw 		: cw_t := "10000011110 1000000110 100000000001100110 0000 0000000 000 000";
	constant bne_cw 		: cw_t := "10000011110 1000000110 100000000001101110 0000 0000000 000 000";
	constant blez_cw 		: cw_t := "10000011110 1000000110 100000000001000110 0000 0000000 000 000";
	constant bgtz_cw 		: cw_t := "10000011110 1000000110 100000000001011110 0000 0000000 000 000";
	constant addi_cw 		: cw_t := "10000011100 1000001000 000000000001000110 1100 0000000 101 100";
	constant addui_cw 		: cw_t := "10000001100 1000001000 000000000000000110 1100 0000000 101 100";
	constant subi_cw 		: cw_t := "10000011100 1000001000 100000000001000110 1100 0000000 101 100";
	constant subui_cw 		: cw_t := "10000001100 1000001000 100000000000000110 1100 0000000 101 100";
	constant andi_cw 		: cw_t := "10000001100 1000001000 000001000110000110 1100 0000000 101 100";
	constant ori_cw 		: cw_t := "10000001100 1000001000 000001110110000110 1100 0000000 101 100";
	constant xori_cw 		: cw_t := "10000001100 1000001000 000000110110000110 1100 0000000 101 100";
	constant beqz_cw 		: cw_t := "10000011110 1000000110 100000000001100110 0000 0000000 000 000";
	constant bnez_cw 		: cw_t := "10000011110 1000000110 100000000001101110 0000 0000000 000 000";
	constant slli_cw 		: cw_t := "10000001100 0010001000 000110000100000110 1100 0000000 101 100";
	constant srli_cw 		: cw_t := "10000001100 0010001000 000100000100000110 1100 0000000 101 100";
	constant srai_cw 		: cw_t := "10000001100 0010001000 001000000100000110 1100 0000000 101 100";
	constant seqi_cw 		: cw_t := "10000011100 1000001000 100000000001000100 1100 0000000 101 100";
	constant snei_cw 		: cw_t := "10000011100 1000001000 100000000001000101 1100 0000000 101 100";
	constant slti_cw 		: cw_t := "10000011100 1000001000 100000000001000001 1100 0000000 101 100";
	constant sgti_cw 		: cw_t := "10000011100 1000001000 100000000001000011 1100 0000000 101 100";
	constant slei_cw 		: cw_t := "10000011100 1000001000 100000000001000000 1100 0000000 101 100";
	constant sgei_cw 		: cw_t := "10000011100 1000001000 100000000001000010 1100 0000000 101 100";
	constant lb_cw			: cw_t := "10000011100 1000001000 000000000001000110 1100 0001100 011 110";
	constant lh_cw	 		: cw_t := "10000011100 1000001000 000000000001000110 1100 0001010 011 110";
	constant lw_cw	 		: cw_t := "10000011100 1000001000 000000000001000110 1100 0001000 011 110";
	constant lbu_cw 		: cw_t := "10000011100 1000001000 000000000001000110 1100 0000100 011 110";
	constant lhu_cw 		: cw_t := "10000011100 1000001000 000000000001000110 1100 0000010 011 110";
	constant sb_cw 			: cw_t := "10000011100 1000000001 000000000001000110 1101 1110001 000 000";
	constant sh_cw 			: cw_t := "10000011100 1000000001 000000000001000110 1101 1100001 000 000";
	constant sw_cw	 		: cw_t := "10000011100 1000000001 000000000001000110 1101 1010001 000 000";
	constant sltui_cw 		: cw_t := "10000011100 1000001000 100000000000000001 1100 0000000 101 100";
	constant sgtui_cw 		: cw_t := "10000011100 1000001000 100000000000000011 1100 0000000 101 100";
	constant sleui_cw 		: cw_t := "10000011100 1000001000 100000000000000000 1100 0000000 101 100";
	constant sgeui_cw 		: cw_t := "10000011100 1000001000 100000000000000010 1100 0000000 101 100";
end package control_words;