library ieee;
use ieee.std_logic_1164.all;

package func_words is
	subtype fw_t is std_logic_vector(62 downto 0);
							   --  ID	        ID/EXE       EXE                E/M     MEM      M/W  WB
	constant nop_fw 	: fw_t	:= "00000001110 001000100000 000110000100111110 0011001 00000000 1011 100";
	constant sll_fw 	: fw_t 	:= "00000001110 001000100010 000110000100111110 0011001 00000000 1011 100";
	constant srl_fw 	: fw_t 	:= "00000001110 001000100010 000100000100111110 0011001 00000000 1011 100";
	constant sra_fw 	: fw_t 	:= "00000001110 001000100010 001000000100111110 0011001 00000000 1011 100";
	constant jr_fw 		: fw_t 	:= "01001101110 100000000001 000000000000110110 0100000 00000000 0000 000";
	constant jalr_fw	: fw_t 	:= "01001101111 100000100101 000000000000110110 0111011 00000001 1011 100";
	constant mult_fw 	: fw_t 	:= "00000001110 010001000010 000000000010111110 0010000 00000000 1000 001";
	constant mfhi_fw 	: fw_t 	:= "00100001110 100000100000 000000000000111110 0011001 00000000 1011 100";
	constant mflo_fw 	: fw_t 	:= "00010001110 100000100000 000000000000111110 0011001 00000000 1011 100";
	constant add_fw 	: fw_t 	:= "00000001110 100000100010 000000000001111110 0011001 00000000 1011 100";
	constant addu_fw 	: fw_t 	:= "00000001110 100000100010 000000000000111110 0011001 00000000 1011 100";
	constant sub_fw 	: fw_t 	:= "00000001110 100000100010 100000000001111110 0011001 00000000 1011 100";
	constant subu_fw 	: fw_t 	:= "00000001110 100000100010 100000000000111110 0011001 00000000 1011 100";
	constant and_fw 	: fw_t 	:= "00000001110 100000100010 000001000110111110 0011001 00000000 1011 100";
	constant or_fw	 	: fw_t 	:= "00000001110 100000100010 000001110110111110 0011001 00000000 1011 100";
	constant xor_fw 	: fw_t 	:= "00000001110 100000100010 000000110110111110 0011001 00000000 1011 100";
	constant seq_fw 	: fw_t 	:= "00000001110 100000100010 100000000001100100 0011001 00000000 1011 100";
	constant sne_fw 	: fw_t 	:= "00000001110 100000100010 100000000001101101 0011001 00000000 1011 100";
	constant slt_fw 	: fw_t 	:= "00000001110 100000100010 100000000001001001 0011001 00000000 1011 100";
	constant sgt_fw 	: fw_t 	:= "00000001110 100000100010 100000000001011011 0011001 00000000 1011 100";
	constant sle_fw 	: fw_t 	:= "00000001110 100000100010 100000000001000000 0011001 00000000 1011 100";
	constant sge_fw 	: fw_t 	:= "00000001110 100000100010 100000000001010010 0011001 00000000 1011 100";
	constant sltu_fw 	: fw_t 	:= "00000001110 100000100010 100000000000001001 0011001 00000000 1011 100";
	constant sgtu_fw 	: fw_t 	:= "00000001110 100000100010 100000000000011011 0011001 00000000 1011 100";
	constant sleu_fw 	: fw_t 	:= "00000001110 100000100010 100000000000000000 0011001 00000000 1011 100";
	constant sgeu_fw 	: fw_t 	:= "00000001110 100000100010 100000000000010010 0011001 00000000 1011 100";
end package func_words;