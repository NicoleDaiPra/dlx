library ieee;
use ieee.std_logic_1164.all;

package func_words is
	subtype fw_t is std_logic_vector(57 downto 0);
							   --  ID	        ID/EXE     EXE                  E/M  MEM     M/W WB
	constant nop_fw 	: fw_t	:= "0000000111000100010000001100001001111100011000000000101100";
	constant sll_fw 	: fw_t 	:= "0000000111000100010000001100001001111100011000000000101100";
	constant srl_fw 	: fw_t 	:= "0000000111000100010000001000001001111100011000000000101100";
	constant sra_fw 	: fw_t 	:= "0000000111000100010000010000001001111100011000000000101100";
	constant jr_fw 		: fw_t 	:= "0100110111010000000000000000000001101100100000000000000000";
	constant jalr_fw	: fw_t 	:= "0100110111110000010010000000000001101100111010000001101100";
	constant mult_fw 	: fw_t 	:= "0000000111001000100000000000000101111100010000000000100001";
	constant mfhi_fw 	: fw_t 	:= "0010000111010000010000000000000001111100011000000000101100";
	constant mflo_fw 	: fw_t 	:= "0001000111010000010000000000000001111100011000000000101100";
	constant add_fw 	: fw_t 	:= "0000000111010000010000000000000011111100011000000000101100";
	constant addu_fw 	: fw_t 	:= "0000000111010000010000000000000001111100011000000000101100";
	constant sub_fw 	: fw_t 	:= "0000000111010000010001000000000011111100011000000000101100";
	constant subu_fw 	: fw_t 	:= "0000000111010000010001000000000001111100011000000000101100";
	constant and_fw 	: fw_t 	:= "0000000111010000010000000010001101111100011000000000101100";
	constant or_fw	 	: fw_t 	:= "0000000111010000010000000011101101111100011000000000101100";
	constant xor_fw 	: fw_t 	:= "0000000111010000010000000001101101111100011000000000101100";
	constant seq_fw 	: fw_t 	:= "0000000111010000010001000000000011111000011000000000101100";
	constant sne_fw 	: fw_t 	:= "0000000111010000010001000000000011111010011000000000101100";
	constant slt_fw 	: fw_t 	:= "0000000111010000010001000000000011110010011000000000101100";
	constant sgt_fw 	: fw_t 	:= "0000000111010000010001000000000011110110011000000000101100";
	constant sle_fw 	: fw_t 	:= "0000000111010000010001000000000011110000011000000000101100";
	constant sge_fw 	: fw_t 	:= "0000000111010000010001000000000011110100011000000000101100";
	constant sltu_fw 	: fw_t 	:= "0000000111010000010001000000000001110010011000000000101100";
	constant sgtu_fw 	: fw_t 	:= "0000000111010000010001000000000001110110011000000000101100";
	constant sleu_fw 	: fw_t 	:= "0000000111010000010001000000000001110000011000000000101100";
	constant sgeu_fw 	: fw_t 	:= "0000000111010000010001000000000001110100011000000000101100";
end package func_words;