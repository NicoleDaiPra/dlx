library ieee;
use ieee.std_logic_1164.all;

package func_words is
	subtype fw_t is std_logic_vector(58 downto 0);
							   --  ID	        ID/EXE     EXE                  E/M  MEM     M/W WB
	constant nop_fw 	: fw_t	:= "00000001110001000100000011000010011111000110000000000101100";
	constant sll_fw 	: fw_t 	:= "00000001110001000100000011000010011111000110000000000101100";
	constant srl_fw 	: fw_t 	:= "00000001110001000100000010000010011111000110000000000101100";
	constant sra_fw 	: fw_t 	:= "00000001110001000100000100000010011111000110000000000101100";
	constant jr_fw 		: fw_t 	:= "01001101110100000000000000000000011011001000000000000000000";
	constant jalr_fw	: fw_t 	:= "01001101111100000100100000000000011011001110100000001101100";
	constant mult_fw 	: fw_t 	:= "00000001110010001000000000000001011111000100000000000100001";
	constant mfhi_fw 	: fw_t 	:= "00100001110100000100000000000000011111000110000000000101100";
	constant mflo_fw 	: fw_t 	:= "00010001110100000100000000000000011111000110000000000101100";
	constant add_fw 	: fw_t 	:= "00000001110100000100000000000000111111000110000000000101100";
	constant addu_fw 	: fw_t 	:= "00000001110100000100000000000000011111000110000000000101100";
	constant sub_fw 	: fw_t 	:= "00000001110100000100010000000000111111000110000000000101100";
	constant subu_fw 	: fw_t 	:= "00000001110100000100010000000000011111000110000000000101100";
	constant and_fw 	: fw_t 	:= "00000001110100000100000000100011011111000110000000000101100";
	constant or_fw	 	: fw_t 	:= "00000001110100000100000000111011011111000110000000000101100";
	constant xor_fw 	: fw_t 	:= "00000001110100000100000000011011011111000110000000000101100";
	constant seq_fw 	: fw_t 	:= "00000001110100000100010000000000110010000110000000000101100";
	constant sne_fw 	: fw_t 	:= "00000001110100000100010000000000110110100110000000000101100";
	constant slt_fw 	: fw_t 	:= "00000001110100000100010000000000100100100110000000000101100";
	constant sgt_fw 	: fw_t 	:= "00000001110100000100010000000000101101100110000000000101100";
	constant sle_fw 	: fw_t 	:= "00000001110100000100010000000000100000000110000000000101100";
	constant sge_fw 	: fw_t 	:= "00000001110100000100010000000000101001000110000000000101100";
	constant sltu_fw 	: fw_t 	:= "00000001110100000100010000000000000100100110000000000101100";
	constant sgtu_fw 	: fw_t 	:= "00000001110100000100010000000000001101100110000000000101100";
	constant sleu_fw 	: fw_t 	:= "00000001110100000100010000000000000000000110000000000101100";
	constant sgeu_fw 	: fw_t 	:= "00000001110100000100010000000000001001000110000000000101100";
end package func_words;