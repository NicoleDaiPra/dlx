
module rf_N32 ( clk, rst, rp1_addr, rp2_addr, wp_addr, wp_en, wp, rp1, rp2, 
        rp1_out_sel, rp2_out_sel, hilo_wr_en, lo_in, hi_in );
  input [4:0] rp1_addr;
  input [4:0] rp2_addr;
  input [4:0] wp_addr;
  input [31:0] wp;
  output [31:0] rp1;
  output [31:0] rp2;
  input [1:0] rp1_out_sel;
  input [1:0] rp2_out_sel;
  input [31:0] lo_in;
  input [31:0] hi_in;
  input clk, rst, wp_en, hilo_wr_en;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n2482, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2623, n2624, n2625, n2626,
         n2627, n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636,
         n2637, n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646,
         n2647, n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656,
         n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666,
         n2667, n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676,
         n2677, n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686,
         n2687, n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696,
         n2697, n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706,
         n2707, n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716,
         n2717, n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726,
         n2727, n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736,
         n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746,
         n2747, n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006,
         n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016,
         n3017, n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026,
         n3027, n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036,
         n3037, n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046,
         n3047, n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066,
         n3067, n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076,
         n3077, n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086,
         n3087, n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096,
         n3097, n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106,
         n3107, n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116,
         n3117, n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126,
         n3127, n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136,
         n3137, n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146,
         n3147, n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156,
         n3157, n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166,
         n3167, n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176,
         n3177, n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186,
         n3187, n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196,
         n3197, n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206,
         n3207, n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216,
         n3217, n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226,
         n3227, n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236,
         n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246,
         n3247, n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256,
         n3257, n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266,
         n3267, n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276,
         n3277, n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286,
         n3287, n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296,
         n3297, n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306,
         n3307, n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316,
         n3317, n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326,
         n3327, n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336,
         n3337, n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346,
         n3347, n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356,
         n3357, n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366,
         n3367, n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376,
         n3377, n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386,
         n3387, n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396,
         n3397, n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406,
         n3407, n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416,
         n3417, n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426,
         n3427, n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436,
         n3437, n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446,
         n3447, n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456,
         n3457, n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466,
         n3467, n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476,
         n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486,
         n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496,
         n3497, n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506,
         n3507, n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516,
         n3517, n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526,
         n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536,
         n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546,
         n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596,
         n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606,
         n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225,
         n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235,
         n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245,
         n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255,
         n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265,
         n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275,
         n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285,
         n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295,
         n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305,
         n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315,
         n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325,
         n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335,
         n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345,
         n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355,
         n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365,
         n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375,
         n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385,
         n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395,
         n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405,
         n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415,
         n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425,
         n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435,
         n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445,
         n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455,
         n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465,
         n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475,
         n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485,
         n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495,
         n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505,
         n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515,
         n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525,
         n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535,
         n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545,
         n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555,
         n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565,
         n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575,
         n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585,
         n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595,
         n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605,
         n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615,
         n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625,
         n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635,
         n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645,
         n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655,
         n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665,
         n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675,
         n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685,
         n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695,
         n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705,
         n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715,
         n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725,
         n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735,
         n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745,
         n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755,
         n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765,
         n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775,
         n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785,
         n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795,
         n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805,
         n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815,
         n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825,
         n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835,
         n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845,
         n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855,
         n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865,
         n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875,
         n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885,
         n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895,
         n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905,
         n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915,
         n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925,
         n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935,
         n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945,
         n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955,
         n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965,
         n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975,
         n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985,
         n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995,
         n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005,
         n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015,
         n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025,
         n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035,
         n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045,
         n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055,
         n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065,
         n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075,
         n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085,
         n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095,
         n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105,
         n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115,
         n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125,
         n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135,
         n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145,
         n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155,
         n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165,
         n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175,
         n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185,
         n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195,
         n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205,
         n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215,
         n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225,
         n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235,
         n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245,
         n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255,
         n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265,
         n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275,
         n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285,
         n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295,
         n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305,
         n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315,
         n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325,
         n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335,
         n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345,
         n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355,
         n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365,
         n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375,
         n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385,
         n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395,
         n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405,
         n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415,
         n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425,
         n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435,
         n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445,
         n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455,
         n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465,
         n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475,
         n2476, n2477, n2478, n2479, n2480, n2481, n2483, n2484, n2548, n2549,
         n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n2620, n2621, n2622, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787;
  wire   [31:0] lo_out;
  wire   [31:0] hi_out;

  DFF_X1 \reg_1/q_reg[0]  ( .D(n3614), .CK(n993), .QN(n1) );
  DFF_X1 \reg_1/q_reg[1]  ( .D(n3613), .CK(n993), .QN(n2) );
  DFF_X1 \reg_1/q_reg[2]  ( .D(n3612), .CK(n993), .QN(n3) );
  DFF_X1 \reg_1/q_reg[3]  ( .D(n3611), .CK(n993), .QN(n4) );
  DFF_X1 \reg_1/q_reg[4]  ( .D(n3610), .CK(n993), .QN(n5) );
  DFF_X1 \reg_1/q_reg[5]  ( .D(n3609), .CK(n993), .QN(n6) );
  DFF_X1 \reg_1/q_reg[6]  ( .D(n3608), .CK(n993), .QN(n7) );
  DFF_X1 \reg_1/q_reg[7]  ( .D(n3607), .CK(n993), .QN(n8) );
  DFF_X1 \reg_1/q_reg[8]  ( .D(n3606), .CK(n993), .QN(n9) );
  DFF_X1 \reg_1/q_reg[9]  ( .D(n3605), .CK(n993), .QN(n10) );
  DFF_X1 \reg_1/q_reg[10]  ( .D(n3604), .CK(n993), .QN(n11) );
  DFF_X1 \reg_1/q_reg[11]  ( .D(n3603), .CK(n993), .QN(n12) );
  DFF_X1 \reg_1/q_reg[12]  ( .D(n3602), .CK(n993), .QN(n13) );
  DFF_X1 \reg_1/q_reg[13]  ( .D(n3601), .CK(n993), .QN(n14) );
  DFF_X1 \reg_1/q_reg[14]  ( .D(n3600), .CK(n993), .QN(n15) );
  DFF_X1 \reg_1/q_reg[15]  ( .D(n3599), .CK(n993), .QN(n16) );
  DFF_X1 \reg_1/q_reg[16]  ( .D(n3598), .CK(n993), .QN(n17) );
  DFF_X1 \reg_1/q_reg[17]  ( .D(n3597), .CK(n993), .QN(n18) );
  DFF_X1 \reg_1/q_reg[18]  ( .D(n3596), .CK(n993), .QN(n19) );
  DFF_X1 \reg_1/q_reg[19]  ( .D(n3595), .CK(n993), .QN(n20) );
  DFF_X1 \reg_1/q_reg[20]  ( .D(n3594), .CK(n993), .QN(n21) );
  DFF_X1 \reg_1/q_reg[21]  ( .D(n3593), .CK(n993), .QN(n22) );
  DFF_X1 \reg_1/q_reg[22]  ( .D(n3592), .CK(n993), .QN(n23) );
  DFF_X1 \reg_1/q_reg[23]  ( .D(n3591), .CK(n993), .QN(n24) );
  DFF_X1 \reg_1/q_reg[24]  ( .D(n3590), .CK(n993), .QN(n25) );
  DFF_X1 \reg_1/q_reg[25]  ( .D(n3589), .CK(n993), .QN(n26) );
  DFF_X1 \reg_1/q_reg[26]  ( .D(n3588), .CK(n993), .QN(n27) );
  DFF_X1 \reg_1/q_reg[27]  ( .D(n3587), .CK(n993), .QN(n28) );
  DFF_X1 \reg_1/q_reg[28]  ( .D(n3586), .CK(n993), .QN(n29) );
  DFF_X1 \reg_1/q_reg[29]  ( .D(n3585), .CK(n993), .QN(n30) );
  DFF_X1 \reg_1/q_reg[30]  ( .D(n3584), .CK(n993), .QN(n31) );
  DFF_X1 \reg_1/q_reg[31]  ( .D(n3583), .CK(n993), .QN(n32) );
  DFF_X1 \reg_2/q_reg[0]  ( .D(n3582), .CK(n993), .QN(n33) );
  DFF_X1 \reg_2/q_reg[1]  ( .D(n3581), .CK(n993), .QN(n34) );
  DFF_X1 \reg_2/q_reg[2]  ( .D(n3580), .CK(n993), .QN(n35) );
  DFF_X1 \reg_2/q_reg[3]  ( .D(n3579), .CK(n993), .QN(n36) );
  DFF_X1 \reg_2/q_reg[4]  ( .D(n3578), .CK(n993), .QN(n37) );
  DFF_X1 \reg_2/q_reg[5]  ( .D(n3577), .CK(n993), .QN(n38) );
  DFF_X1 \reg_2/q_reg[6]  ( .D(n3576), .CK(n993), .QN(n39) );
  DFF_X1 \reg_2/q_reg[7]  ( .D(n3575), .CK(n993), .QN(n40) );
  DFF_X1 \reg_2/q_reg[8]  ( .D(n3574), .CK(n993), .QN(n41) );
  DFF_X1 \reg_2/q_reg[9]  ( .D(n3573), .CK(n993), .QN(n42) );
  DFF_X1 \reg_2/q_reg[10]  ( .D(n3572), .CK(n993), .QN(n43) );
  DFF_X1 \reg_2/q_reg[11]  ( .D(n3571), .CK(n993), .QN(n44) );
  DFF_X1 \reg_2/q_reg[12]  ( .D(n3570), .CK(n993), .QN(n45) );
  DFF_X1 \reg_2/q_reg[13]  ( .D(n3569), .CK(n993), .QN(n46) );
  DFF_X1 \reg_2/q_reg[14]  ( .D(n3568), .CK(n993), .QN(n47) );
  DFF_X1 \reg_2/q_reg[15]  ( .D(n3567), .CK(n993), .QN(n48) );
  DFF_X1 \reg_2/q_reg[16]  ( .D(n3566), .CK(n993), .QN(n49) );
  DFF_X1 \reg_2/q_reg[17]  ( .D(n3565), .CK(n993), .QN(n50) );
  DFF_X1 \reg_2/q_reg[18]  ( .D(n3564), .CK(n993), .QN(n51) );
  DFF_X1 \reg_2/q_reg[19]  ( .D(n3563), .CK(n993), .QN(n52) );
  DFF_X1 \reg_2/q_reg[20]  ( .D(n3562), .CK(n993), .QN(n53) );
  DFF_X1 \reg_2/q_reg[21]  ( .D(n3561), .CK(n993), .QN(n54) );
  DFF_X1 \reg_2/q_reg[22]  ( .D(n3560), .CK(n993), .QN(n55) );
  DFF_X1 \reg_2/q_reg[23]  ( .D(n3559), .CK(n993), .QN(n56) );
  DFF_X1 \reg_2/q_reg[24]  ( .D(n3558), .CK(n993), .QN(n57) );
  DFF_X1 \reg_2/q_reg[25]  ( .D(n3557), .CK(n993), .QN(n58) );
  DFF_X1 \reg_2/q_reg[26]  ( .D(n3556), .CK(n993), .QN(n59) );
  DFF_X1 \reg_2/q_reg[27]  ( .D(n3555), .CK(n993), .QN(n60) );
  DFF_X1 \reg_2/q_reg[28]  ( .D(n3554), .CK(n993), .QN(n61) );
  DFF_X1 \reg_2/q_reg[29]  ( .D(n3553), .CK(n993), .QN(n62) );
  DFF_X1 \reg_2/q_reg[30]  ( .D(n3552), .CK(n993), .QN(n63) );
  DFF_X1 \reg_2/q_reg[31]  ( .D(n3551), .CK(n993), .QN(n64) );
  DFF_X1 \reg_3/q_reg[0]  ( .D(n3550), .CK(n993), .QN(n65) );
  DFF_X1 \reg_3/q_reg[1]  ( .D(n3549), .CK(n993), .QN(n66) );
  DFF_X1 \reg_3/q_reg[2]  ( .D(n3548), .CK(n993), .QN(n67) );
  DFF_X1 \reg_3/q_reg[3]  ( .D(n3547), .CK(n993), .QN(n68) );
  DFF_X1 \reg_3/q_reg[4]  ( .D(n3546), .CK(n993), .QN(n69) );
  DFF_X1 \reg_3/q_reg[5]  ( .D(n3545), .CK(n993), .QN(n70) );
  DFF_X1 \reg_3/q_reg[6]  ( .D(n3544), .CK(n993), .QN(n71) );
  DFF_X1 \reg_3/q_reg[7]  ( .D(n3543), .CK(n993), .QN(n72) );
  DFF_X1 \reg_3/q_reg[8]  ( .D(n3542), .CK(n993), .QN(n73) );
  DFF_X1 \reg_3/q_reg[9]  ( .D(n3541), .CK(n993), .QN(n74) );
  DFF_X1 \reg_3/q_reg[10]  ( .D(n3540), .CK(n993), .QN(n75) );
  DFF_X1 \reg_3/q_reg[11]  ( .D(n3539), .CK(n993), .QN(n76) );
  DFF_X1 \reg_3/q_reg[12]  ( .D(n3538), .CK(n993), .QN(n77) );
  DFF_X1 \reg_3/q_reg[13]  ( .D(n3537), .CK(n993), .QN(n78) );
  DFF_X1 \reg_3/q_reg[14]  ( .D(n3536), .CK(n993), .QN(n79) );
  DFF_X1 \reg_3/q_reg[15]  ( .D(n3535), .CK(n993), .QN(n80) );
  DFF_X1 \reg_3/q_reg[16]  ( .D(n3534), .CK(n993), .QN(n81) );
  DFF_X1 \reg_3/q_reg[17]  ( .D(n3533), .CK(n993), .QN(n82) );
  DFF_X1 \reg_3/q_reg[18]  ( .D(n3532), .CK(n993), .QN(n83) );
  DFF_X1 \reg_3/q_reg[19]  ( .D(n3531), .CK(n993), .QN(n84) );
  DFF_X1 \reg_3/q_reg[20]  ( .D(n3530), .CK(n993), .QN(n85) );
  DFF_X1 \reg_3/q_reg[21]  ( .D(n3529), .CK(n993), .QN(n86) );
  DFF_X1 \reg_3/q_reg[22]  ( .D(n3528), .CK(n993), .QN(n87) );
  DFF_X1 \reg_3/q_reg[23]  ( .D(n3527), .CK(n993), .QN(n88) );
  DFF_X1 \reg_3/q_reg[24]  ( .D(n3526), .CK(n993), .QN(n89) );
  DFF_X1 \reg_3/q_reg[25]  ( .D(n3525), .CK(n993), .QN(n90) );
  DFF_X1 \reg_3/q_reg[26]  ( .D(n3524), .CK(n993), .QN(n91) );
  DFF_X1 \reg_3/q_reg[27]  ( .D(n3523), .CK(n993), .QN(n92) );
  DFF_X1 \reg_3/q_reg[28]  ( .D(n3522), .CK(n993), .QN(n93) );
  DFF_X1 \reg_3/q_reg[29]  ( .D(n3521), .CK(n993), .QN(n94) );
  DFF_X1 \reg_3/q_reg[30]  ( .D(n3520), .CK(n993), .QN(n95) );
  DFF_X1 \reg_3/q_reg[31]  ( .D(n3519), .CK(n993), .QN(n96) );
  DFF_X1 \reg_4/q_reg[0]  ( .D(n3518), .CK(n993), .QN(n97) );
  DFF_X1 \reg_4/q_reg[1]  ( .D(n3517), .CK(n993), .QN(n98) );
  DFF_X1 \reg_4/q_reg[2]  ( .D(n3516), .CK(n993), .QN(n99) );
  DFF_X1 \reg_4/q_reg[3]  ( .D(n3515), .CK(n993), .QN(n100) );
  DFF_X1 \reg_4/q_reg[4]  ( .D(n3514), .CK(n993), .QN(n101) );
  DFF_X1 \reg_4/q_reg[5]  ( .D(n3513), .CK(n993), .QN(n102) );
  DFF_X1 \reg_4/q_reg[6]  ( .D(n3512), .CK(n993), .QN(n103) );
  DFF_X1 \reg_4/q_reg[7]  ( .D(n3511), .CK(n993), .QN(n104) );
  DFF_X1 \reg_4/q_reg[8]  ( .D(n3510), .CK(n993), .QN(n105) );
  DFF_X1 \reg_4/q_reg[9]  ( .D(n3509), .CK(n993), .QN(n106) );
  DFF_X1 \reg_4/q_reg[10]  ( .D(n3508), .CK(n993), .QN(n107) );
  DFF_X1 \reg_4/q_reg[11]  ( .D(n3507), .CK(n993), .QN(n108) );
  DFF_X1 \reg_4/q_reg[12]  ( .D(n3506), .CK(n993), .QN(n109) );
  DFF_X1 \reg_4/q_reg[13]  ( .D(n3505), .CK(n993), .QN(n110) );
  DFF_X1 \reg_4/q_reg[14]  ( .D(n3504), .CK(n993), .QN(n111) );
  DFF_X1 \reg_4/q_reg[15]  ( .D(n3503), .CK(n993), .QN(n112) );
  DFF_X1 \reg_4/q_reg[16]  ( .D(n3502), .CK(n993), .QN(n113) );
  DFF_X1 \reg_4/q_reg[17]  ( .D(n3501), .CK(n993), .QN(n114) );
  DFF_X1 \reg_4/q_reg[18]  ( .D(n3500), .CK(n993), .QN(n115) );
  DFF_X1 \reg_4/q_reg[19]  ( .D(n3499), .CK(n993), .QN(n116) );
  DFF_X1 \reg_4/q_reg[20]  ( .D(n3498), .CK(n993), .QN(n117) );
  DFF_X1 \reg_4/q_reg[21]  ( .D(n3497), .CK(n993), .QN(n118) );
  DFF_X1 \reg_4/q_reg[22]  ( .D(n3496), .CK(n993), .QN(n119) );
  DFF_X1 \reg_4/q_reg[23]  ( .D(n3495), .CK(n993), .QN(n120) );
  DFF_X1 \reg_4/q_reg[24]  ( .D(n3494), .CK(n993), .QN(n121) );
  DFF_X1 \reg_4/q_reg[25]  ( .D(n3493), .CK(n993), .QN(n122) );
  DFF_X1 \reg_4/q_reg[26]  ( .D(n3492), .CK(n993), .QN(n123) );
  DFF_X1 \reg_4/q_reg[27]  ( .D(n3491), .CK(n993), .QN(n124) );
  DFF_X1 \reg_4/q_reg[28]  ( .D(n3490), .CK(n993), .QN(n125) );
  DFF_X1 \reg_4/q_reg[29]  ( .D(n3489), .CK(n993), .QN(n126) );
  DFF_X1 \reg_4/q_reg[30]  ( .D(n3488), .CK(n993), .QN(n127) );
  DFF_X1 \reg_4/q_reg[31]  ( .D(n3487), .CK(n993), .QN(n128) );
  DFF_X1 \reg_5/q_reg[0]  ( .D(n3486), .CK(n993), .QN(n129) );
  DFF_X1 \reg_5/q_reg[1]  ( .D(n3485), .CK(n993), .QN(n130) );
  DFF_X1 \reg_5/q_reg[2]  ( .D(n3484), .CK(n993), .QN(n131) );
  DFF_X1 \reg_5/q_reg[3]  ( .D(n3483), .CK(n993), .QN(n132) );
  DFF_X1 \reg_5/q_reg[4]  ( .D(n3482), .CK(n993), .QN(n133) );
  DFF_X1 \reg_5/q_reg[5]  ( .D(n3481), .CK(n993), .QN(n134) );
  DFF_X1 \reg_5/q_reg[6]  ( .D(n3480), .CK(n993), .QN(n135) );
  DFF_X1 \reg_5/q_reg[7]  ( .D(n3479), .CK(n993), .QN(n136) );
  DFF_X1 \reg_5/q_reg[8]  ( .D(n3478), .CK(n993), .QN(n137) );
  DFF_X1 \reg_5/q_reg[9]  ( .D(n3477), .CK(n993), .QN(n138) );
  DFF_X1 \reg_5/q_reg[10]  ( .D(n3476), .CK(n993), .QN(n139) );
  DFF_X1 \reg_5/q_reg[11]  ( .D(n3475), .CK(n993), .QN(n140) );
  DFF_X1 \reg_5/q_reg[12]  ( .D(n3474), .CK(n993), .QN(n141) );
  DFF_X1 \reg_5/q_reg[13]  ( .D(n3473), .CK(n993), .QN(n142) );
  DFF_X1 \reg_5/q_reg[14]  ( .D(n3472), .CK(n993), .QN(n143) );
  DFF_X1 \reg_5/q_reg[15]  ( .D(n3471), .CK(n993), .QN(n144) );
  DFF_X1 \reg_5/q_reg[16]  ( .D(n3470), .CK(n993), .QN(n145) );
  DFF_X1 \reg_5/q_reg[17]  ( .D(n3469), .CK(n993), .QN(n146) );
  DFF_X1 \reg_5/q_reg[18]  ( .D(n3468), .CK(n993), .QN(n147) );
  DFF_X1 \reg_5/q_reg[19]  ( .D(n3467), .CK(n993), .QN(n148) );
  DFF_X1 \reg_5/q_reg[20]  ( .D(n3466), .CK(n993), .QN(n149) );
  DFF_X1 \reg_5/q_reg[21]  ( .D(n3465), .CK(n993), .QN(n150) );
  DFF_X1 \reg_5/q_reg[22]  ( .D(n3464), .CK(n993), .QN(n151) );
  DFF_X1 \reg_5/q_reg[23]  ( .D(n3463), .CK(n993), .QN(n152) );
  DFF_X1 \reg_5/q_reg[24]  ( .D(n3462), .CK(n993), .QN(n153) );
  DFF_X1 \reg_5/q_reg[25]  ( .D(n3461), .CK(n993), .QN(n154) );
  DFF_X1 \reg_5/q_reg[26]  ( .D(n3460), .CK(n993), .QN(n155) );
  DFF_X1 \reg_5/q_reg[27]  ( .D(n3459), .CK(n993), .QN(n156) );
  DFF_X1 \reg_5/q_reg[28]  ( .D(n3458), .CK(n993), .QN(n157) );
  DFF_X1 \reg_5/q_reg[29]  ( .D(n3457), .CK(n993), .QN(n158) );
  DFF_X1 \reg_5/q_reg[30]  ( .D(n3456), .CK(n993), .QN(n159) );
  DFF_X1 \reg_5/q_reg[31]  ( .D(n3455), .CK(n993), .QN(n160) );
  DFF_X1 \reg_6/q_reg[0]  ( .D(n3454), .CK(n993), .QN(n161) );
  DFF_X1 \reg_6/q_reg[1]  ( .D(n3453), .CK(n993), .QN(n162) );
  DFF_X1 \reg_6/q_reg[2]  ( .D(n3452), .CK(n993), .QN(n163) );
  DFF_X1 \reg_6/q_reg[3]  ( .D(n3451), .CK(n993), .QN(n164) );
  DFF_X1 \reg_6/q_reg[4]  ( .D(n3450), .CK(n993), .QN(n165) );
  DFF_X1 \reg_6/q_reg[5]  ( .D(n3449), .CK(n993), .QN(n166) );
  DFF_X1 \reg_6/q_reg[6]  ( .D(n3448), .CK(n993), .QN(n167) );
  DFF_X1 \reg_6/q_reg[7]  ( .D(n3447), .CK(n993), .QN(n168) );
  DFF_X1 \reg_6/q_reg[8]  ( .D(n3446), .CK(n993), .QN(n169) );
  DFF_X1 \reg_6/q_reg[9]  ( .D(n3445), .CK(n993), .QN(n170) );
  DFF_X1 \reg_6/q_reg[10]  ( .D(n3444), .CK(n993), .QN(n171) );
  DFF_X1 \reg_6/q_reg[11]  ( .D(n3443), .CK(n993), .QN(n172) );
  DFF_X1 \reg_6/q_reg[12]  ( .D(n3442), .CK(n993), .QN(n173) );
  DFF_X1 \reg_6/q_reg[13]  ( .D(n3441), .CK(n993), .QN(n174) );
  DFF_X1 \reg_6/q_reg[14]  ( .D(n3440), .CK(n993), .QN(n175) );
  DFF_X1 \reg_6/q_reg[15]  ( .D(n3439), .CK(n993), .QN(n176) );
  DFF_X1 \reg_6/q_reg[16]  ( .D(n3438), .CK(n993), .QN(n177) );
  DFF_X1 \reg_6/q_reg[17]  ( .D(n3437), .CK(n993), .QN(n178) );
  DFF_X1 \reg_6/q_reg[18]  ( .D(n3436), .CK(n993), .QN(n179) );
  DFF_X1 \reg_6/q_reg[19]  ( .D(n3435), .CK(n993), .QN(n180) );
  DFF_X1 \reg_6/q_reg[20]  ( .D(n3434), .CK(n993), .QN(n181) );
  DFF_X1 \reg_6/q_reg[21]  ( .D(n3433), .CK(n993), .QN(n182) );
  DFF_X1 \reg_6/q_reg[22]  ( .D(n3432), .CK(n993), .QN(n183) );
  DFF_X1 \reg_6/q_reg[23]  ( .D(n3431), .CK(n993), .QN(n184) );
  DFF_X1 \reg_6/q_reg[24]  ( .D(n3430), .CK(n993), .QN(n185) );
  DFF_X1 \reg_6/q_reg[25]  ( .D(n3429), .CK(n993), .QN(n186) );
  DFF_X1 \reg_6/q_reg[26]  ( .D(n3428), .CK(n993), .QN(n187) );
  DFF_X1 \reg_6/q_reg[27]  ( .D(n3427), .CK(n993), .QN(n188) );
  DFF_X1 \reg_6/q_reg[28]  ( .D(n3426), .CK(n993), .QN(n189) );
  DFF_X1 \reg_6/q_reg[29]  ( .D(n3425), .CK(n993), .QN(n190) );
  DFF_X1 \reg_6/q_reg[30]  ( .D(n3424), .CK(n993), .QN(n191) );
  DFF_X1 \reg_6/q_reg[31]  ( .D(n3423), .CK(n993), .QN(n192) );
  DFF_X1 \reg_7/q_reg[0]  ( .D(n3422), .CK(n993), .QN(n193) );
  DFF_X1 \reg_7/q_reg[1]  ( .D(n3421), .CK(n993), .QN(n194) );
  DFF_X1 \reg_7/q_reg[2]  ( .D(n3420), .CK(n993), .QN(n195) );
  DFF_X1 \reg_7/q_reg[3]  ( .D(n3419), .CK(n993), .QN(n196) );
  DFF_X1 \reg_7/q_reg[4]  ( .D(n3418), .CK(n993), .QN(n197) );
  DFF_X1 \reg_7/q_reg[5]  ( .D(n3417), .CK(n993), .QN(n198) );
  DFF_X1 \reg_7/q_reg[6]  ( .D(n3416), .CK(n993), .QN(n199) );
  DFF_X1 \reg_7/q_reg[7]  ( .D(n3415), .CK(n993), .QN(n200) );
  DFF_X1 \reg_7/q_reg[8]  ( .D(n3414), .CK(n993), .QN(n201) );
  DFF_X1 \reg_7/q_reg[9]  ( .D(n3413), .CK(n993), .QN(n202) );
  DFF_X1 \reg_7/q_reg[10]  ( .D(n3412), .CK(n993), .QN(n203) );
  DFF_X1 \reg_7/q_reg[11]  ( .D(n3411), .CK(n993), .QN(n204) );
  DFF_X1 \reg_7/q_reg[12]  ( .D(n3410), .CK(n993), .QN(n205) );
  DFF_X1 \reg_7/q_reg[13]  ( .D(n3409), .CK(n993), .QN(n206) );
  DFF_X1 \reg_7/q_reg[14]  ( .D(n3408), .CK(n993), .QN(n207) );
  DFF_X1 \reg_7/q_reg[15]  ( .D(n3407), .CK(n993), .QN(n208) );
  DFF_X1 \reg_7/q_reg[16]  ( .D(n3406), .CK(n993), .QN(n209) );
  DFF_X1 \reg_7/q_reg[17]  ( .D(n3405), .CK(n993), .QN(n210) );
  DFF_X1 \reg_7/q_reg[18]  ( .D(n3404), .CK(n993), .QN(n211) );
  DFF_X1 \reg_7/q_reg[19]  ( .D(n3403), .CK(n993), .QN(n212) );
  DFF_X1 \reg_7/q_reg[20]  ( .D(n3402), .CK(n993), .QN(n213) );
  DFF_X1 \reg_7/q_reg[21]  ( .D(n3401), .CK(n993), .QN(n214) );
  DFF_X1 \reg_7/q_reg[22]  ( .D(n3400), .CK(n993), .QN(n215) );
  DFF_X1 \reg_7/q_reg[23]  ( .D(n3399), .CK(n993), .QN(n216) );
  DFF_X1 \reg_7/q_reg[24]  ( .D(n3398), .CK(n993), .QN(n217) );
  DFF_X1 \reg_7/q_reg[25]  ( .D(n3397), .CK(n993), .QN(n218) );
  DFF_X1 \reg_7/q_reg[26]  ( .D(n3396), .CK(n993), .QN(n219) );
  DFF_X1 \reg_7/q_reg[27]  ( .D(n3395), .CK(n993), .QN(n220) );
  DFF_X1 \reg_7/q_reg[28]  ( .D(n3394), .CK(n993), .QN(n221) );
  DFF_X1 \reg_7/q_reg[29]  ( .D(n3393), .CK(n993), .QN(n222) );
  DFF_X1 \reg_7/q_reg[30]  ( .D(n3392), .CK(n993), .QN(n223) );
  DFF_X1 \reg_7/q_reg[31]  ( .D(n3391), .CK(n993), .QN(n224) );
  DFF_X1 \reg_8/q_reg[0]  ( .D(n3390), .CK(n993), .QN(n225) );
  DFF_X1 \reg_8/q_reg[1]  ( .D(n3389), .CK(n993), .QN(n226) );
  DFF_X1 \reg_8/q_reg[2]  ( .D(n3388), .CK(n993), .QN(n227) );
  DFF_X1 \reg_8/q_reg[3]  ( .D(n3387), .CK(n993), .QN(n228) );
  DFF_X1 \reg_8/q_reg[4]  ( .D(n3386), .CK(n993), .QN(n229) );
  DFF_X1 \reg_8/q_reg[5]  ( .D(n3385), .CK(n993), .QN(n230) );
  DFF_X1 \reg_8/q_reg[6]  ( .D(n3384), .CK(n993), .QN(n231) );
  DFF_X1 \reg_8/q_reg[7]  ( .D(n3383), .CK(n993), .QN(n232) );
  DFF_X1 \reg_8/q_reg[8]  ( .D(n3382), .CK(n993), .QN(n233) );
  DFF_X1 \reg_8/q_reg[9]  ( .D(n3381), .CK(n993), .QN(n234) );
  DFF_X1 \reg_8/q_reg[10]  ( .D(n3380), .CK(n993), .QN(n235) );
  DFF_X1 \reg_8/q_reg[11]  ( .D(n3379), .CK(n993), .QN(n236) );
  DFF_X1 \reg_8/q_reg[12]  ( .D(n3378), .CK(n993), .QN(n237) );
  DFF_X1 \reg_8/q_reg[13]  ( .D(n3377), .CK(n993), .QN(n238) );
  DFF_X1 \reg_8/q_reg[14]  ( .D(n3376), .CK(n993), .QN(n239) );
  DFF_X1 \reg_8/q_reg[15]  ( .D(n3375), .CK(n993), .QN(n240) );
  DFF_X1 \reg_8/q_reg[16]  ( .D(n3374), .CK(n993), .QN(n241) );
  DFF_X1 \reg_8/q_reg[17]  ( .D(n3373), .CK(n993), .QN(n242) );
  DFF_X1 \reg_8/q_reg[18]  ( .D(n3372), .CK(n993), .QN(n243) );
  DFF_X1 \reg_8/q_reg[19]  ( .D(n3371), .CK(n993), .QN(n244) );
  DFF_X1 \reg_8/q_reg[20]  ( .D(n3370), .CK(n993), .QN(n245) );
  DFF_X1 \reg_8/q_reg[21]  ( .D(n3369), .CK(n993), .QN(n246) );
  DFF_X1 \reg_8/q_reg[22]  ( .D(n3368), .CK(n993), .QN(n247) );
  DFF_X1 \reg_8/q_reg[23]  ( .D(n3367), .CK(n993), .QN(n248) );
  DFF_X1 \reg_8/q_reg[24]  ( .D(n3366), .CK(n993), .QN(n249) );
  DFF_X1 \reg_8/q_reg[25]  ( .D(n3365), .CK(n993), .QN(n250) );
  DFF_X1 \reg_8/q_reg[26]  ( .D(n3364), .CK(n993), .QN(n251) );
  DFF_X1 \reg_8/q_reg[27]  ( .D(n3363), .CK(n993), .QN(n252) );
  DFF_X1 \reg_8/q_reg[28]  ( .D(n3362), .CK(n993), .QN(n253) );
  DFF_X1 \reg_8/q_reg[29]  ( .D(n3361), .CK(n993), .QN(n254) );
  DFF_X1 \reg_8/q_reg[30]  ( .D(n3360), .CK(n993), .QN(n255) );
  DFF_X1 \reg_8/q_reg[31]  ( .D(n3359), .CK(n993), .QN(n256) );
  DFF_X1 \reg_9/q_reg[0]  ( .D(n3358), .CK(n993), .QN(n257) );
  DFF_X1 \reg_9/q_reg[1]  ( .D(n3357), .CK(n993), .QN(n258) );
  DFF_X1 \reg_9/q_reg[2]  ( .D(n3356), .CK(n993), .QN(n259) );
  DFF_X1 \reg_9/q_reg[3]  ( .D(n3355), .CK(n993), .QN(n260) );
  DFF_X1 \reg_9/q_reg[4]  ( .D(n3354), .CK(n993), .QN(n261) );
  DFF_X1 \reg_9/q_reg[5]  ( .D(n3353), .CK(n993), .QN(n262) );
  DFF_X1 \reg_9/q_reg[6]  ( .D(n3352), .CK(n993), .QN(n263) );
  DFF_X1 \reg_9/q_reg[7]  ( .D(n3351), .CK(n993), .QN(n264) );
  DFF_X1 \reg_9/q_reg[8]  ( .D(n3350), .CK(n993), .QN(n265) );
  DFF_X1 \reg_9/q_reg[9]  ( .D(n3349), .CK(n993), .QN(n266) );
  DFF_X1 \reg_9/q_reg[10]  ( .D(n3348), .CK(n993), .QN(n267) );
  DFF_X1 \reg_9/q_reg[11]  ( .D(n3347), .CK(n993), .QN(n268) );
  DFF_X1 \reg_9/q_reg[12]  ( .D(n3346), .CK(n993), .QN(n269) );
  DFF_X1 \reg_9/q_reg[13]  ( .D(n3345), .CK(n993), .QN(n270) );
  DFF_X1 \reg_9/q_reg[14]  ( .D(n3344), .CK(n993), .QN(n271) );
  DFF_X1 \reg_9/q_reg[15]  ( .D(n3343), .CK(n993), .QN(n272) );
  DFF_X1 \reg_9/q_reg[16]  ( .D(n3342), .CK(n993), .QN(n273) );
  DFF_X1 \reg_9/q_reg[17]  ( .D(n3341), .CK(n993), .QN(n274) );
  DFF_X1 \reg_9/q_reg[18]  ( .D(n3340), .CK(n993), .QN(n275) );
  DFF_X1 \reg_9/q_reg[19]  ( .D(n3339), .CK(n993), .QN(n276) );
  DFF_X1 \reg_9/q_reg[20]  ( .D(n3338), .CK(n993), .QN(n277) );
  DFF_X1 \reg_9/q_reg[21]  ( .D(n3337), .CK(n993), .QN(n278) );
  DFF_X1 \reg_9/q_reg[22]  ( .D(n3336), .CK(n993), .QN(n279) );
  DFF_X1 \reg_9/q_reg[23]  ( .D(n3335), .CK(n993), .QN(n280) );
  DFF_X1 \reg_9/q_reg[24]  ( .D(n3334), .CK(n993), .QN(n281) );
  DFF_X1 \reg_9/q_reg[25]  ( .D(n3333), .CK(n993), .QN(n282) );
  DFF_X1 \reg_9/q_reg[26]  ( .D(n3332), .CK(n993), .QN(n283) );
  DFF_X1 \reg_9/q_reg[27]  ( .D(n3331), .CK(n993), .QN(n284) );
  DFF_X1 \reg_9/q_reg[28]  ( .D(n3330), .CK(n993), .QN(n285) );
  DFF_X1 \reg_9/q_reg[29]  ( .D(n3329), .CK(n993), .QN(n286) );
  DFF_X1 \reg_9/q_reg[30]  ( .D(n3328), .CK(n993), .QN(n287) );
  DFF_X1 \reg_9/q_reg[31]  ( .D(n3327), .CK(n993), .QN(n288) );
  DFF_X1 \reg_10/q_reg[0]  ( .D(n3326), .CK(n993), .QN(n289) );
  DFF_X1 \reg_10/q_reg[1]  ( .D(n3325), .CK(n993), .QN(n290) );
  DFF_X1 \reg_10/q_reg[2]  ( .D(n3324), .CK(n993), .QN(n291) );
  DFF_X1 \reg_10/q_reg[3]  ( .D(n3323), .CK(n993), .QN(n292) );
  DFF_X1 \reg_10/q_reg[4]  ( .D(n3322), .CK(n993), .QN(n293) );
  DFF_X1 \reg_10/q_reg[5]  ( .D(n3321), .CK(n993), .QN(n294) );
  DFF_X1 \reg_10/q_reg[6]  ( .D(n3320), .CK(n993), .QN(n295) );
  DFF_X1 \reg_10/q_reg[7]  ( .D(n3319), .CK(n993), .QN(n296) );
  DFF_X1 \reg_10/q_reg[8]  ( .D(n3318), .CK(n993), .QN(n297) );
  DFF_X1 \reg_10/q_reg[9]  ( .D(n3317), .CK(n993), .QN(n298) );
  DFF_X1 \reg_10/q_reg[10]  ( .D(n3316), .CK(n993), .QN(n299) );
  DFF_X1 \reg_10/q_reg[11]  ( .D(n3315), .CK(n993), .QN(n300) );
  DFF_X1 \reg_10/q_reg[12]  ( .D(n3314), .CK(n993), .QN(n301) );
  DFF_X1 \reg_10/q_reg[13]  ( .D(n3313), .CK(n993), .QN(n302) );
  DFF_X1 \reg_10/q_reg[14]  ( .D(n3312), .CK(n993), .QN(n303) );
  DFF_X1 \reg_10/q_reg[15]  ( .D(n3311), .CK(n993), .QN(n304) );
  DFF_X1 \reg_10/q_reg[16]  ( .D(n3310), .CK(n993), .QN(n305) );
  DFF_X1 \reg_10/q_reg[17]  ( .D(n3309), .CK(n993), .QN(n306) );
  DFF_X1 \reg_10/q_reg[18]  ( .D(n3308), .CK(n993), .QN(n307) );
  DFF_X1 \reg_10/q_reg[19]  ( .D(n3307), .CK(n993), .QN(n308) );
  DFF_X1 \reg_10/q_reg[20]  ( .D(n3306), .CK(n993), .QN(n309) );
  DFF_X1 \reg_10/q_reg[21]  ( .D(n3305), .CK(n993), .QN(n310) );
  DFF_X1 \reg_10/q_reg[22]  ( .D(n3304), .CK(n993), .QN(n311) );
  DFF_X1 \reg_10/q_reg[23]  ( .D(n3303), .CK(n993), .QN(n312) );
  DFF_X1 \reg_10/q_reg[24]  ( .D(n3302), .CK(n993), .QN(n313) );
  DFF_X1 \reg_10/q_reg[25]  ( .D(n3301), .CK(n993), .QN(n314) );
  DFF_X1 \reg_10/q_reg[26]  ( .D(n3300), .CK(n993), .QN(n315) );
  DFF_X1 \reg_10/q_reg[27]  ( .D(n3299), .CK(n993), .QN(n316) );
  DFF_X1 \reg_10/q_reg[28]  ( .D(n3298), .CK(n993), .QN(n317) );
  DFF_X1 \reg_10/q_reg[29]  ( .D(n3297), .CK(n993), .QN(n318) );
  DFF_X1 \reg_10/q_reg[30]  ( .D(n3296), .CK(n993), .QN(n319) );
  DFF_X1 \reg_10/q_reg[31]  ( .D(n3295), .CK(n993), .QN(n320) );
  DFF_X1 \reg_11/q_reg[0]  ( .D(n3294), .CK(n993), .QN(n321) );
  DFF_X1 \reg_11/q_reg[1]  ( .D(n3293), .CK(n993), .QN(n322) );
  DFF_X1 \reg_11/q_reg[2]  ( .D(n3292), .CK(n993), .QN(n323) );
  DFF_X1 \reg_11/q_reg[3]  ( .D(n3291), .CK(n993), .QN(n324) );
  DFF_X1 \reg_11/q_reg[4]  ( .D(n3290), .CK(n993), .QN(n325) );
  DFF_X1 \reg_11/q_reg[5]  ( .D(n3289), .CK(n993), .QN(n326) );
  DFF_X1 \reg_11/q_reg[6]  ( .D(n3288), .CK(n993), .QN(n327) );
  DFF_X1 \reg_11/q_reg[7]  ( .D(n3287), .CK(n993), .QN(n328) );
  DFF_X1 \reg_11/q_reg[8]  ( .D(n3286), .CK(n993), .QN(n329) );
  DFF_X1 \reg_11/q_reg[9]  ( .D(n3285), .CK(n993), .QN(n330) );
  DFF_X1 \reg_11/q_reg[10]  ( .D(n3284), .CK(n993), .QN(n331) );
  DFF_X1 \reg_11/q_reg[11]  ( .D(n3283), .CK(n993), .QN(n332) );
  DFF_X1 \reg_11/q_reg[12]  ( .D(n3282), .CK(n993), .QN(n333) );
  DFF_X1 \reg_11/q_reg[13]  ( .D(n3281), .CK(n993), .QN(n334) );
  DFF_X1 \reg_11/q_reg[14]  ( .D(n3280), .CK(n993), .QN(n335) );
  DFF_X1 \reg_11/q_reg[15]  ( .D(n3279), .CK(n993), .QN(n336) );
  DFF_X1 \reg_11/q_reg[16]  ( .D(n3278), .CK(n993), .QN(n337) );
  DFF_X1 \reg_11/q_reg[17]  ( .D(n3277), .CK(n993), .QN(n338) );
  DFF_X1 \reg_11/q_reg[18]  ( .D(n3276), .CK(n993), .QN(n339) );
  DFF_X1 \reg_11/q_reg[19]  ( .D(n3275), .CK(n993), .QN(n340) );
  DFF_X1 \reg_11/q_reg[20]  ( .D(n3274), .CK(n993), .QN(n341) );
  DFF_X1 \reg_11/q_reg[21]  ( .D(n3273), .CK(n993), .QN(n342) );
  DFF_X1 \reg_11/q_reg[22]  ( .D(n3272), .CK(n993), .QN(n343) );
  DFF_X1 \reg_11/q_reg[23]  ( .D(n3271), .CK(n993), .QN(n344) );
  DFF_X1 \reg_11/q_reg[24]  ( .D(n3270), .CK(n993), .QN(n345) );
  DFF_X1 \reg_11/q_reg[25]  ( .D(n3269), .CK(n993), .QN(n346) );
  DFF_X1 \reg_11/q_reg[26]  ( .D(n3268), .CK(n993), .QN(n347) );
  DFF_X1 \reg_11/q_reg[27]  ( .D(n3267), .CK(n993), .QN(n348) );
  DFF_X1 \reg_11/q_reg[28]  ( .D(n3266), .CK(n993), .QN(n349) );
  DFF_X1 \reg_11/q_reg[29]  ( .D(n3265), .CK(n993), .QN(n350) );
  DFF_X1 \reg_11/q_reg[30]  ( .D(n3264), .CK(n993), .QN(n351) );
  DFF_X1 \reg_11/q_reg[31]  ( .D(n3263), .CK(n993), .QN(n352) );
  DFF_X1 \reg_12/q_reg[0]  ( .D(n3262), .CK(n993), .QN(n353) );
  DFF_X1 \reg_12/q_reg[1]  ( .D(n3261), .CK(n993), .QN(n354) );
  DFF_X1 \reg_12/q_reg[2]  ( .D(n3260), .CK(n993), .QN(n355) );
  DFF_X1 \reg_12/q_reg[3]  ( .D(n3259), .CK(n993), .QN(n356) );
  DFF_X1 \reg_12/q_reg[4]  ( .D(n3258), .CK(n993), .QN(n357) );
  DFF_X1 \reg_12/q_reg[5]  ( .D(n3257), .CK(n993), .QN(n358) );
  DFF_X1 \reg_12/q_reg[6]  ( .D(n3256), .CK(n993), .QN(n359) );
  DFF_X1 \reg_12/q_reg[7]  ( .D(n3255), .CK(n993), .QN(n360) );
  DFF_X1 \reg_12/q_reg[8]  ( .D(n3254), .CK(n993), .QN(n361) );
  DFF_X1 \reg_12/q_reg[9]  ( .D(n3253), .CK(n993), .QN(n362) );
  DFF_X1 \reg_12/q_reg[10]  ( .D(n3252), .CK(n993), .QN(n363) );
  DFF_X1 \reg_12/q_reg[11]  ( .D(n3251), .CK(n993), .QN(n364) );
  DFF_X1 \reg_12/q_reg[12]  ( .D(n3250), .CK(n993), .QN(n365) );
  DFF_X1 \reg_12/q_reg[13]  ( .D(n3249), .CK(n993), .QN(n366) );
  DFF_X1 \reg_12/q_reg[14]  ( .D(n3248), .CK(n993), .QN(n367) );
  DFF_X1 \reg_12/q_reg[15]  ( .D(n3247), .CK(n993), .QN(n368) );
  DFF_X1 \reg_12/q_reg[16]  ( .D(n3246), .CK(n993), .QN(n369) );
  DFF_X1 \reg_12/q_reg[17]  ( .D(n3245), .CK(n993), .QN(n370) );
  DFF_X1 \reg_12/q_reg[18]  ( .D(n3244), .CK(n993), .QN(n371) );
  DFF_X1 \reg_12/q_reg[19]  ( .D(n3243), .CK(n993), .QN(n372) );
  DFF_X1 \reg_12/q_reg[20]  ( .D(n3242), .CK(n993), .QN(n373) );
  DFF_X1 \reg_12/q_reg[21]  ( .D(n3241), .CK(n993), .QN(n374) );
  DFF_X1 \reg_12/q_reg[22]  ( .D(n3240), .CK(n993), .QN(n375) );
  DFF_X1 \reg_12/q_reg[23]  ( .D(n3239), .CK(n993), .QN(n376) );
  DFF_X1 \reg_12/q_reg[24]  ( .D(n3238), .CK(n993), .QN(n377) );
  DFF_X1 \reg_12/q_reg[25]  ( .D(n3237), .CK(n993), .QN(n378) );
  DFF_X1 \reg_12/q_reg[26]  ( .D(n3236), .CK(n993), .QN(n379) );
  DFF_X1 \reg_12/q_reg[27]  ( .D(n3235), .CK(n993), .QN(n380) );
  DFF_X1 \reg_12/q_reg[28]  ( .D(n3234), .CK(n993), .QN(n381) );
  DFF_X1 \reg_12/q_reg[29]  ( .D(n3233), .CK(n993), .QN(n382) );
  DFF_X1 \reg_12/q_reg[30]  ( .D(n3232), .CK(n993), .QN(n383) );
  DFF_X1 \reg_12/q_reg[31]  ( .D(n3231), .CK(n993), .QN(n384) );
  DFF_X1 \reg_13/q_reg[0]  ( .D(n3230), .CK(n993), .QN(n385) );
  DFF_X1 \reg_13/q_reg[1]  ( .D(n3229), .CK(n993), .QN(n386) );
  DFF_X1 \reg_13/q_reg[2]  ( .D(n3228), .CK(n993), .QN(n387) );
  DFF_X1 \reg_13/q_reg[3]  ( .D(n3227), .CK(n993), .QN(n388) );
  DFF_X1 \reg_13/q_reg[4]  ( .D(n3226), .CK(n993), .QN(n389) );
  DFF_X1 \reg_13/q_reg[5]  ( .D(n3225), .CK(n993), .QN(n390) );
  DFF_X1 \reg_13/q_reg[6]  ( .D(n3224), .CK(n993), .QN(n391) );
  DFF_X1 \reg_13/q_reg[7]  ( .D(n3223), .CK(n993), .QN(n392) );
  DFF_X1 \reg_13/q_reg[8]  ( .D(n3222), .CK(n993), .QN(n393) );
  DFF_X1 \reg_13/q_reg[9]  ( .D(n3221), .CK(n993), .QN(n394) );
  DFF_X1 \reg_13/q_reg[10]  ( .D(n3220), .CK(n993), .QN(n395) );
  DFF_X1 \reg_13/q_reg[11]  ( .D(n3219), .CK(n993), .QN(n396) );
  DFF_X1 \reg_13/q_reg[12]  ( .D(n3218), .CK(n993), .QN(n397) );
  DFF_X1 \reg_13/q_reg[13]  ( .D(n3217), .CK(n993), .QN(n398) );
  DFF_X1 \reg_13/q_reg[14]  ( .D(n3216), .CK(n993), .QN(n399) );
  DFF_X1 \reg_13/q_reg[15]  ( .D(n3215), .CK(n993), .QN(n400) );
  DFF_X1 \reg_13/q_reg[16]  ( .D(n3214), .CK(n993), .QN(n401) );
  DFF_X1 \reg_13/q_reg[17]  ( .D(n3213), .CK(n993), .QN(n402) );
  DFF_X1 \reg_13/q_reg[18]  ( .D(n3212), .CK(n993), .QN(n403) );
  DFF_X1 \reg_13/q_reg[19]  ( .D(n3211), .CK(n993), .QN(n404) );
  DFF_X1 \reg_13/q_reg[20]  ( .D(n3210), .CK(n993), .QN(n405) );
  DFF_X1 \reg_13/q_reg[21]  ( .D(n3209), .CK(n993), .QN(n406) );
  DFF_X1 \reg_13/q_reg[22]  ( .D(n3208), .CK(n993), .QN(n407) );
  DFF_X1 \reg_13/q_reg[23]  ( .D(n3207), .CK(n993), .QN(n408) );
  DFF_X1 \reg_13/q_reg[24]  ( .D(n3206), .CK(n993), .QN(n409) );
  DFF_X1 \reg_13/q_reg[25]  ( .D(n3205), .CK(n993), .QN(n410) );
  DFF_X1 \reg_13/q_reg[26]  ( .D(n3204), .CK(n993), .QN(n411) );
  DFF_X1 \reg_13/q_reg[27]  ( .D(n3203), .CK(n993), .QN(n412) );
  DFF_X1 \reg_13/q_reg[28]  ( .D(n3202), .CK(n993), .QN(n413) );
  DFF_X1 \reg_13/q_reg[29]  ( .D(n3201), .CK(n993), .QN(n414) );
  DFF_X1 \reg_13/q_reg[30]  ( .D(n3200), .CK(n993), .QN(n415) );
  DFF_X1 \reg_13/q_reg[31]  ( .D(n3199), .CK(n993), .QN(n416) );
  DFF_X1 \reg_14/q_reg[0]  ( .D(n3198), .CK(n993), .QN(n417) );
  DFF_X1 \reg_14/q_reg[1]  ( .D(n3197), .CK(n993), .QN(n418) );
  DFF_X1 \reg_14/q_reg[2]  ( .D(n3196), .CK(n993), .QN(n419) );
  DFF_X1 \reg_14/q_reg[3]  ( .D(n3195), .CK(n993), .QN(n420) );
  DFF_X1 \reg_14/q_reg[4]  ( .D(n3194), .CK(n993), .QN(n421) );
  DFF_X1 \reg_14/q_reg[5]  ( .D(n3193), .CK(n993), .QN(n422) );
  DFF_X1 \reg_14/q_reg[6]  ( .D(n3192), .CK(n993), .QN(n423) );
  DFF_X1 \reg_14/q_reg[7]  ( .D(n3191), .CK(n993), .QN(n424) );
  DFF_X1 \reg_14/q_reg[8]  ( .D(n3190), .CK(n993), .QN(n425) );
  DFF_X1 \reg_14/q_reg[9]  ( .D(n3189), .CK(n993), .QN(n426) );
  DFF_X1 \reg_14/q_reg[10]  ( .D(n3188), .CK(n993), .QN(n427) );
  DFF_X1 \reg_14/q_reg[11]  ( .D(n3187), .CK(n993), .QN(n428) );
  DFF_X1 \reg_14/q_reg[12]  ( .D(n3186), .CK(n993), .QN(n429) );
  DFF_X1 \reg_14/q_reg[13]  ( .D(n3185), .CK(n993), .QN(n430) );
  DFF_X1 \reg_14/q_reg[14]  ( .D(n3184), .CK(n993), .QN(n431) );
  DFF_X1 \reg_14/q_reg[15]  ( .D(n3183), .CK(n993), .QN(n432) );
  DFF_X1 \reg_14/q_reg[16]  ( .D(n3182), .CK(n993), .QN(n433) );
  DFF_X1 \reg_14/q_reg[17]  ( .D(n3181), .CK(n993), .QN(n434) );
  DFF_X1 \reg_14/q_reg[18]  ( .D(n3180), .CK(n993), .QN(n435) );
  DFF_X1 \reg_14/q_reg[19]  ( .D(n3179), .CK(n993), .QN(n436) );
  DFF_X1 \reg_14/q_reg[20]  ( .D(n3178), .CK(n993), .QN(n437) );
  DFF_X1 \reg_14/q_reg[21]  ( .D(n3177), .CK(n993), .QN(n438) );
  DFF_X1 \reg_14/q_reg[22]  ( .D(n3176), .CK(n993), .QN(n439) );
  DFF_X1 \reg_14/q_reg[23]  ( .D(n3175), .CK(n993), .QN(n440) );
  DFF_X1 \reg_14/q_reg[24]  ( .D(n3174), .CK(n993), .QN(n441) );
  DFF_X1 \reg_14/q_reg[25]  ( .D(n3173), .CK(n993), .QN(n442) );
  DFF_X1 \reg_14/q_reg[26]  ( .D(n3172), .CK(n993), .QN(n443) );
  DFF_X1 \reg_14/q_reg[27]  ( .D(n3171), .CK(n993), .QN(n444) );
  DFF_X1 \reg_14/q_reg[28]  ( .D(n3170), .CK(n993), .QN(n445) );
  DFF_X1 \reg_14/q_reg[29]  ( .D(n3169), .CK(n993), .QN(n446) );
  DFF_X1 \reg_14/q_reg[30]  ( .D(n3168), .CK(n993), .QN(n447) );
  DFF_X1 \reg_14/q_reg[31]  ( .D(n3167), .CK(n993), .QN(n448) );
  DFF_X1 \reg_15/q_reg[0]  ( .D(n3166), .CK(n993), .QN(n449) );
  DFF_X1 \reg_15/q_reg[1]  ( .D(n3165), .CK(n993), .QN(n450) );
  DFF_X1 \reg_15/q_reg[2]  ( .D(n3164), .CK(n993), .QN(n451) );
  DFF_X1 \reg_15/q_reg[3]  ( .D(n3163), .CK(n993), .QN(n452) );
  DFF_X1 \reg_15/q_reg[4]  ( .D(n3162), .CK(n993), .QN(n453) );
  DFF_X1 \reg_15/q_reg[5]  ( .D(n3161), .CK(n993), .QN(n454) );
  DFF_X1 \reg_15/q_reg[6]  ( .D(n3160), .CK(n993), .QN(n455) );
  DFF_X1 \reg_15/q_reg[7]  ( .D(n3159), .CK(n993), .QN(n456) );
  DFF_X1 \reg_15/q_reg[8]  ( .D(n3158), .CK(n993), .QN(n457) );
  DFF_X1 \reg_15/q_reg[9]  ( .D(n3157), .CK(n993), .QN(n458) );
  DFF_X1 \reg_15/q_reg[10]  ( .D(n3156), .CK(n993), .QN(n459) );
  DFF_X1 \reg_15/q_reg[11]  ( .D(n3155), .CK(n993), .QN(n460) );
  DFF_X1 \reg_15/q_reg[12]  ( .D(n3154), .CK(n993), .QN(n461) );
  DFF_X1 \reg_15/q_reg[13]  ( .D(n3153), .CK(n993), .QN(n462) );
  DFF_X1 \reg_15/q_reg[14]  ( .D(n3152), .CK(n993), .QN(n463) );
  DFF_X1 \reg_15/q_reg[15]  ( .D(n3151), .CK(n993), .QN(n464) );
  DFF_X1 \reg_15/q_reg[16]  ( .D(n3150), .CK(n993), .QN(n465) );
  DFF_X1 \reg_15/q_reg[17]  ( .D(n3149), .CK(n993), .QN(n466) );
  DFF_X1 \reg_15/q_reg[18]  ( .D(n3148), .CK(n993), .QN(n467) );
  DFF_X1 \reg_15/q_reg[19]  ( .D(n3147), .CK(n993), .QN(n468) );
  DFF_X1 \reg_15/q_reg[20]  ( .D(n3146), .CK(n993), .QN(n469) );
  DFF_X1 \reg_15/q_reg[21]  ( .D(n3145), .CK(n993), .QN(n470) );
  DFF_X1 \reg_15/q_reg[22]  ( .D(n3144), .CK(n993), .QN(n471) );
  DFF_X1 \reg_15/q_reg[23]  ( .D(n3143), .CK(n993), .QN(n472) );
  DFF_X1 \reg_15/q_reg[24]  ( .D(n3142), .CK(n993), .QN(n473) );
  DFF_X1 \reg_15/q_reg[25]  ( .D(n3141), .CK(n993), .QN(n474) );
  DFF_X1 \reg_15/q_reg[26]  ( .D(n3140), .CK(n993), .QN(n475) );
  DFF_X1 \reg_15/q_reg[27]  ( .D(n3139), .CK(n993), .QN(n476) );
  DFF_X1 \reg_15/q_reg[28]  ( .D(n3138), .CK(n993), .QN(n477) );
  DFF_X1 \reg_15/q_reg[29]  ( .D(n3137), .CK(n993), .QN(n478) );
  DFF_X1 \reg_15/q_reg[30]  ( .D(n3136), .CK(n993), .QN(n479) );
  DFF_X1 \reg_15/q_reg[31]  ( .D(n3135), .CK(n993), .QN(n480) );
  DFF_X1 \reg_16/q_reg[0]  ( .D(n3134), .CK(n993), .QN(n481) );
  DFF_X1 \reg_16/q_reg[1]  ( .D(n3133), .CK(n993), .QN(n482) );
  DFF_X1 \reg_16/q_reg[2]  ( .D(n3132), .CK(n993), .QN(n483) );
  DFF_X1 \reg_16/q_reg[3]  ( .D(n3131), .CK(n993), .QN(n484) );
  DFF_X1 \reg_16/q_reg[4]  ( .D(n3130), .CK(n993), .QN(n485) );
  DFF_X1 \reg_16/q_reg[5]  ( .D(n3129), .CK(n993), .QN(n486) );
  DFF_X1 \reg_16/q_reg[6]  ( .D(n3128), .CK(n993), .QN(n487) );
  DFF_X1 \reg_16/q_reg[7]  ( .D(n3127), .CK(n993), .QN(n488) );
  DFF_X1 \reg_16/q_reg[8]  ( .D(n3126), .CK(n993), .QN(n489) );
  DFF_X1 \reg_16/q_reg[9]  ( .D(n3125), .CK(n993), .QN(n490) );
  DFF_X1 \reg_16/q_reg[10]  ( .D(n3124), .CK(n993), .QN(n491) );
  DFF_X1 \reg_16/q_reg[11]  ( .D(n3123), .CK(n993), .QN(n492) );
  DFF_X1 \reg_16/q_reg[12]  ( .D(n3122), .CK(n993), .QN(n493) );
  DFF_X1 \reg_16/q_reg[13]  ( .D(n3121), .CK(n993), .QN(n494) );
  DFF_X1 \reg_16/q_reg[14]  ( .D(n3120), .CK(n993), .QN(n495) );
  DFF_X1 \reg_16/q_reg[15]  ( .D(n3119), .CK(n993), .QN(n496) );
  DFF_X1 \reg_16/q_reg[16]  ( .D(n3118), .CK(n993), .QN(n497) );
  DFF_X1 \reg_16/q_reg[17]  ( .D(n3117), .CK(n993), .QN(n498) );
  DFF_X1 \reg_16/q_reg[18]  ( .D(n3116), .CK(n993), .QN(n499) );
  DFF_X1 \reg_16/q_reg[19]  ( .D(n3115), .CK(n993), .QN(n500) );
  DFF_X1 \reg_16/q_reg[20]  ( .D(n3114), .CK(n993), .QN(n501) );
  DFF_X1 \reg_16/q_reg[21]  ( .D(n3113), .CK(n993), .QN(n502) );
  DFF_X1 \reg_16/q_reg[22]  ( .D(n3112), .CK(n993), .QN(n503) );
  DFF_X1 \reg_16/q_reg[23]  ( .D(n3111), .CK(n993), .QN(n504) );
  DFF_X1 \reg_16/q_reg[24]  ( .D(n3110), .CK(n993), .QN(n505) );
  DFF_X1 \reg_16/q_reg[25]  ( .D(n3109), .CK(n993), .QN(n506) );
  DFF_X1 \reg_16/q_reg[26]  ( .D(n3108), .CK(n993), .QN(n507) );
  DFF_X1 \reg_16/q_reg[27]  ( .D(n3107), .CK(n993), .QN(n508) );
  DFF_X1 \reg_16/q_reg[28]  ( .D(n3106), .CK(n993), .QN(n509) );
  DFF_X1 \reg_16/q_reg[29]  ( .D(n3105), .CK(n993), .QN(n510) );
  DFF_X1 \reg_16/q_reg[30]  ( .D(n3104), .CK(n993), .QN(n511) );
  DFF_X1 \reg_16/q_reg[31]  ( .D(n3103), .CK(n993), .QN(n512) );
  DFF_X1 \reg_17/q_reg[0]  ( .D(n3102), .CK(n993), .QN(n513) );
  DFF_X1 \reg_17/q_reg[1]  ( .D(n3101), .CK(n993), .QN(n514) );
  DFF_X1 \reg_17/q_reg[2]  ( .D(n3100), .CK(n993), .QN(n515) );
  DFF_X1 \reg_17/q_reg[3]  ( .D(n3099), .CK(n993), .QN(n516) );
  DFF_X1 \reg_17/q_reg[4]  ( .D(n3098), .CK(n993), .QN(n517) );
  DFF_X1 \reg_17/q_reg[5]  ( .D(n3097), .CK(n993), .QN(n518) );
  DFF_X1 \reg_17/q_reg[6]  ( .D(n3096), .CK(n993), .QN(n519) );
  DFF_X1 \reg_17/q_reg[7]  ( .D(n3095), .CK(n993), .QN(n520) );
  DFF_X1 \reg_17/q_reg[8]  ( .D(n3094), .CK(n993), .QN(n521) );
  DFF_X1 \reg_17/q_reg[9]  ( .D(n3093), .CK(n993), .QN(n522) );
  DFF_X1 \reg_17/q_reg[10]  ( .D(n3092), .CK(n993), .QN(n523) );
  DFF_X1 \reg_17/q_reg[11]  ( .D(n3091), .CK(n993), .QN(n524) );
  DFF_X1 \reg_17/q_reg[12]  ( .D(n3090), .CK(n993), .QN(n525) );
  DFF_X1 \reg_17/q_reg[13]  ( .D(n3089), .CK(n993), .QN(n526) );
  DFF_X1 \reg_17/q_reg[14]  ( .D(n3088), .CK(n993), .QN(n527) );
  DFF_X1 \reg_17/q_reg[15]  ( .D(n3087), .CK(n993), .QN(n528) );
  DFF_X1 \reg_17/q_reg[16]  ( .D(n3086), .CK(n993), .QN(n529) );
  DFF_X1 \reg_17/q_reg[17]  ( .D(n3085), .CK(n993), .QN(n530) );
  DFF_X1 \reg_17/q_reg[18]  ( .D(n3084), .CK(n993), .QN(n531) );
  DFF_X1 \reg_17/q_reg[19]  ( .D(n3083), .CK(n993), .QN(n532) );
  DFF_X1 \reg_17/q_reg[20]  ( .D(n3082), .CK(n993), .QN(n533) );
  DFF_X1 \reg_17/q_reg[21]  ( .D(n3081), .CK(n993), .QN(n534) );
  DFF_X1 \reg_17/q_reg[22]  ( .D(n3080), .CK(n993), .QN(n535) );
  DFF_X1 \reg_17/q_reg[23]  ( .D(n3079), .CK(n993), .QN(n536) );
  DFF_X1 \reg_17/q_reg[24]  ( .D(n3078), .CK(n993), .QN(n537) );
  DFF_X1 \reg_17/q_reg[25]  ( .D(n3077), .CK(n993), .QN(n538) );
  DFF_X1 \reg_17/q_reg[26]  ( .D(n3076), .CK(n993), .QN(n539) );
  DFF_X1 \reg_17/q_reg[27]  ( .D(n3075), .CK(n993), .QN(n540) );
  DFF_X1 \reg_17/q_reg[28]  ( .D(n3074), .CK(n993), .QN(n541) );
  DFF_X1 \reg_17/q_reg[29]  ( .D(n3073), .CK(n993), .QN(n542) );
  DFF_X1 \reg_17/q_reg[30]  ( .D(n3072), .CK(n993), .QN(n543) );
  DFF_X1 \reg_17/q_reg[31]  ( .D(n3071), .CK(n993), .QN(n544) );
  DFF_X1 \reg_18/q_reg[0]  ( .D(n3070), .CK(n993), .QN(n545) );
  DFF_X1 \reg_18/q_reg[1]  ( .D(n3069), .CK(n993), .QN(n546) );
  DFF_X1 \reg_18/q_reg[2]  ( .D(n3068), .CK(n993), .QN(n547) );
  DFF_X1 \reg_18/q_reg[3]  ( .D(n3067), .CK(n993), .QN(n548) );
  DFF_X1 \reg_18/q_reg[4]  ( .D(n3066), .CK(n993), .QN(n549) );
  DFF_X1 \reg_18/q_reg[5]  ( .D(n3065), .CK(n993), .QN(n550) );
  DFF_X1 \reg_18/q_reg[6]  ( .D(n3064), .CK(n993), .QN(n551) );
  DFF_X1 \reg_18/q_reg[7]  ( .D(n3063), .CK(n993), .QN(n552) );
  DFF_X1 \reg_18/q_reg[8]  ( .D(n3062), .CK(n993), .QN(n553) );
  DFF_X1 \reg_18/q_reg[9]  ( .D(n3061), .CK(n993), .QN(n554) );
  DFF_X1 \reg_18/q_reg[10]  ( .D(n3060), .CK(n993), .QN(n555) );
  DFF_X1 \reg_18/q_reg[11]  ( .D(n3059), .CK(n993), .QN(n556) );
  DFF_X1 \reg_18/q_reg[12]  ( .D(n3058), .CK(n993), .QN(n557) );
  DFF_X1 \reg_18/q_reg[13]  ( .D(n3057), .CK(n993), .QN(n558) );
  DFF_X1 \reg_18/q_reg[14]  ( .D(n3056), .CK(n993), .QN(n559) );
  DFF_X1 \reg_18/q_reg[15]  ( .D(n3055), .CK(n993), .QN(n560) );
  DFF_X1 \reg_18/q_reg[16]  ( .D(n3054), .CK(n993), .QN(n561) );
  DFF_X1 \reg_18/q_reg[17]  ( .D(n3053), .CK(n993), .QN(n562) );
  DFF_X1 \reg_18/q_reg[18]  ( .D(n3052), .CK(n993), .QN(n563) );
  DFF_X1 \reg_18/q_reg[19]  ( .D(n3051), .CK(n993), .QN(n564) );
  DFF_X1 \reg_18/q_reg[20]  ( .D(n3050), .CK(n993), .QN(n565) );
  DFF_X1 \reg_18/q_reg[21]  ( .D(n3049), .CK(n993), .QN(n566) );
  DFF_X1 \reg_18/q_reg[22]  ( .D(n3048), .CK(n993), .QN(n567) );
  DFF_X1 \reg_18/q_reg[23]  ( .D(n3047), .CK(n993), .QN(n568) );
  DFF_X1 \reg_18/q_reg[24]  ( .D(n3046), .CK(n993), .QN(n569) );
  DFF_X1 \reg_18/q_reg[25]  ( .D(n3045), .CK(n993), .QN(n570) );
  DFF_X1 \reg_18/q_reg[26]  ( .D(n3044), .CK(n993), .QN(n571) );
  DFF_X1 \reg_18/q_reg[27]  ( .D(n3043), .CK(n993), .QN(n572) );
  DFF_X1 \reg_18/q_reg[28]  ( .D(n3042), .CK(n993), .QN(n573) );
  DFF_X1 \reg_18/q_reg[29]  ( .D(n3041), .CK(n993), .QN(n574) );
  DFF_X1 \reg_18/q_reg[30]  ( .D(n3040), .CK(n993), .QN(n575) );
  DFF_X1 \reg_18/q_reg[31]  ( .D(n3039), .CK(n993), .QN(n576) );
  DFF_X1 \reg_19/q_reg[0]  ( .D(n3038), .CK(n993), .QN(n577) );
  DFF_X1 \reg_19/q_reg[1]  ( .D(n3037), .CK(n993), .QN(n578) );
  DFF_X1 \reg_19/q_reg[2]  ( .D(n3036), .CK(n993), .QN(n579) );
  DFF_X1 \reg_19/q_reg[3]  ( .D(n3035), .CK(n993), .QN(n580) );
  DFF_X1 \reg_19/q_reg[4]  ( .D(n3034), .CK(n993), .QN(n581) );
  DFF_X1 \reg_19/q_reg[5]  ( .D(n3033), .CK(n993), .QN(n582) );
  DFF_X1 \reg_19/q_reg[6]  ( .D(n3032), .CK(n993), .QN(n583) );
  DFF_X1 \reg_19/q_reg[7]  ( .D(n3031), .CK(n993), .QN(n584) );
  DFF_X1 \reg_19/q_reg[8]  ( .D(n3030), .CK(n993), .QN(n585) );
  DFF_X1 \reg_19/q_reg[9]  ( .D(n3029), .CK(n993), .QN(n586) );
  DFF_X1 \reg_19/q_reg[10]  ( .D(n3028), .CK(n993), .QN(n587) );
  DFF_X1 \reg_19/q_reg[11]  ( .D(n3027), .CK(n993), .QN(n588) );
  DFF_X1 \reg_19/q_reg[12]  ( .D(n3026), .CK(n993), .QN(n589) );
  DFF_X1 \reg_19/q_reg[13]  ( .D(n3025), .CK(n993), .QN(n590) );
  DFF_X1 \reg_19/q_reg[14]  ( .D(n3024), .CK(n993), .QN(n591) );
  DFF_X1 \reg_19/q_reg[15]  ( .D(n3023), .CK(n993), .QN(n592) );
  DFF_X1 \reg_19/q_reg[16]  ( .D(n3022), .CK(n993), .QN(n593) );
  DFF_X1 \reg_19/q_reg[17]  ( .D(n3021), .CK(n993), .QN(n594) );
  DFF_X1 \reg_19/q_reg[18]  ( .D(n3020), .CK(n993), .QN(n595) );
  DFF_X1 \reg_19/q_reg[19]  ( .D(n3019), .CK(n993), .QN(n596) );
  DFF_X1 \reg_19/q_reg[20]  ( .D(n3018), .CK(n993), .QN(n597) );
  DFF_X1 \reg_19/q_reg[21]  ( .D(n3017), .CK(n993), .QN(n598) );
  DFF_X1 \reg_19/q_reg[22]  ( .D(n3016), .CK(n993), .QN(n599) );
  DFF_X1 \reg_19/q_reg[23]  ( .D(n3015), .CK(n993), .QN(n600) );
  DFF_X1 \reg_19/q_reg[24]  ( .D(n3014), .CK(n993), .QN(n601) );
  DFF_X1 \reg_19/q_reg[25]  ( .D(n3013), .CK(n993), .QN(n602) );
  DFF_X1 \reg_19/q_reg[26]  ( .D(n3012), .CK(n993), .QN(n603) );
  DFF_X1 \reg_19/q_reg[27]  ( .D(n3011), .CK(n993), .QN(n604) );
  DFF_X1 \reg_19/q_reg[28]  ( .D(n3010), .CK(n993), .QN(n605) );
  DFF_X1 \reg_19/q_reg[29]  ( .D(n3009), .CK(n993), .QN(n606) );
  DFF_X1 \reg_19/q_reg[30]  ( .D(n3008), .CK(n993), .QN(n607) );
  DFF_X1 \reg_19/q_reg[31]  ( .D(n3007), .CK(n993), .QN(n608) );
  DFF_X1 \reg_20/q_reg[0]  ( .D(n3006), .CK(n993), .QN(n609) );
  DFF_X1 \reg_20/q_reg[1]  ( .D(n3005), .CK(n993), .QN(n610) );
  DFF_X1 \reg_20/q_reg[2]  ( .D(n3004), .CK(n993), .QN(n611) );
  DFF_X1 \reg_20/q_reg[3]  ( .D(n3003), .CK(n993), .QN(n612) );
  DFF_X1 \reg_20/q_reg[4]  ( .D(n3002), .CK(n993), .QN(n613) );
  DFF_X1 \reg_20/q_reg[5]  ( .D(n3001), .CK(n993), .QN(n614) );
  DFF_X1 \reg_20/q_reg[6]  ( .D(n3000), .CK(n993), .QN(n615) );
  DFF_X1 \reg_20/q_reg[7]  ( .D(n2999), .CK(n993), .QN(n616) );
  DFF_X1 \reg_20/q_reg[8]  ( .D(n2998), .CK(n993), .QN(n617) );
  DFF_X1 \reg_20/q_reg[9]  ( .D(n2997), .CK(n993), .QN(n618) );
  DFF_X1 \reg_20/q_reg[10]  ( .D(n2996), .CK(n993), .QN(n619) );
  DFF_X1 \reg_20/q_reg[11]  ( .D(n2995), .CK(n993), .QN(n620) );
  DFF_X1 \reg_20/q_reg[12]  ( .D(n2994), .CK(n993), .QN(n621) );
  DFF_X1 \reg_20/q_reg[13]  ( .D(n2993), .CK(n993), .QN(n622) );
  DFF_X1 \reg_20/q_reg[14]  ( .D(n2992), .CK(n993), .QN(n623) );
  DFF_X1 \reg_20/q_reg[15]  ( .D(n2991), .CK(n993), .QN(n624) );
  DFF_X1 \reg_20/q_reg[16]  ( .D(n2990), .CK(n993), .QN(n625) );
  DFF_X1 \reg_20/q_reg[17]  ( .D(n2989), .CK(n993), .QN(n626) );
  DFF_X1 \reg_20/q_reg[18]  ( .D(n2988), .CK(n993), .QN(n627) );
  DFF_X1 \reg_20/q_reg[19]  ( .D(n2987), .CK(n993), .QN(n628) );
  DFF_X1 \reg_20/q_reg[20]  ( .D(n2986), .CK(n993), .QN(n629) );
  DFF_X1 \reg_20/q_reg[21]  ( .D(n2985), .CK(n993), .QN(n630) );
  DFF_X1 \reg_20/q_reg[22]  ( .D(n2984), .CK(n993), .QN(n631) );
  DFF_X1 \reg_20/q_reg[23]  ( .D(n2983), .CK(n993), .QN(n632) );
  DFF_X1 \reg_20/q_reg[24]  ( .D(n2982), .CK(n993), .QN(n633) );
  DFF_X1 \reg_20/q_reg[25]  ( .D(n2981), .CK(n993), .QN(n634) );
  DFF_X1 \reg_20/q_reg[26]  ( .D(n2980), .CK(n993), .QN(n635) );
  DFF_X1 \reg_20/q_reg[27]  ( .D(n2979), .CK(n993), .QN(n636) );
  DFF_X1 \reg_20/q_reg[28]  ( .D(n2978), .CK(n993), .QN(n637) );
  DFF_X1 \reg_20/q_reg[29]  ( .D(n2977), .CK(n993), .QN(n638) );
  DFF_X1 \reg_20/q_reg[30]  ( .D(n2976), .CK(n993), .QN(n639) );
  DFF_X1 \reg_20/q_reg[31]  ( .D(n2975), .CK(n993), .QN(n640) );
  DFF_X1 \reg_21/q_reg[0]  ( .D(n2974), .CK(n993), .QN(n641) );
  DFF_X1 \reg_21/q_reg[1]  ( .D(n2973), .CK(n993), .QN(n642) );
  DFF_X1 \reg_21/q_reg[2]  ( .D(n2972), .CK(n993), .QN(n643) );
  DFF_X1 \reg_21/q_reg[3]  ( .D(n2971), .CK(n993), .QN(n644) );
  DFF_X1 \reg_21/q_reg[4]  ( .D(n2970), .CK(n993), .QN(n645) );
  DFF_X1 \reg_21/q_reg[5]  ( .D(n2969), .CK(n993), .QN(n646) );
  DFF_X1 \reg_21/q_reg[6]  ( .D(n2968), .CK(n993), .QN(n647) );
  DFF_X1 \reg_21/q_reg[7]  ( .D(n2967), .CK(n993), .QN(n648) );
  DFF_X1 \reg_21/q_reg[8]  ( .D(n2966), .CK(n993), .QN(n649) );
  DFF_X1 \reg_21/q_reg[9]  ( .D(n2965), .CK(n993), .QN(n650) );
  DFF_X1 \reg_21/q_reg[10]  ( .D(n2964), .CK(n993), .QN(n651) );
  DFF_X1 \reg_21/q_reg[11]  ( .D(n2963), .CK(n993), .QN(n652) );
  DFF_X1 \reg_21/q_reg[12]  ( .D(n2962), .CK(n993), .QN(n653) );
  DFF_X1 \reg_21/q_reg[13]  ( .D(n2961), .CK(n993), .QN(n654) );
  DFF_X1 \reg_21/q_reg[14]  ( .D(n2960), .CK(n993), .QN(n655) );
  DFF_X1 \reg_21/q_reg[15]  ( .D(n2959), .CK(n993), .QN(n656) );
  DFF_X1 \reg_21/q_reg[16]  ( .D(n2958), .CK(n993), .QN(n657) );
  DFF_X1 \reg_21/q_reg[17]  ( .D(n2957), .CK(n993), .QN(n658) );
  DFF_X1 \reg_21/q_reg[18]  ( .D(n2956), .CK(n993), .QN(n659) );
  DFF_X1 \reg_21/q_reg[19]  ( .D(n2955), .CK(n993), .QN(n660) );
  DFF_X1 \reg_21/q_reg[20]  ( .D(n2954), .CK(n993), .QN(n661) );
  DFF_X1 \reg_21/q_reg[21]  ( .D(n2953), .CK(n993), .QN(n662) );
  DFF_X1 \reg_21/q_reg[22]  ( .D(n2952), .CK(n993), .QN(n663) );
  DFF_X1 \reg_21/q_reg[23]  ( .D(n2951), .CK(n993), .QN(n664) );
  DFF_X1 \reg_21/q_reg[24]  ( .D(n2950), .CK(n993), .QN(n665) );
  DFF_X1 \reg_21/q_reg[25]  ( .D(n2949), .CK(n993), .QN(n666) );
  DFF_X1 \reg_21/q_reg[26]  ( .D(n2948), .CK(n993), .QN(n667) );
  DFF_X1 \reg_21/q_reg[27]  ( .D(n2947), .CK(n993), .QN(n668) );
  DFF_X1 \reg_21/q_reg[28]  ( .D(n2946), .CK(n993), .QN(n669) );
  DFF_X1 \reg_21/q_reg[29]  ( .D(n2945), .CK(n993), .QN(n670) );
  DFF_X1 \reg_21/q_reg[30]  ( .D(n2944), .CK(n993), .QN(n671) );
  DFF_X1 \reg_21/q_reg[31]  ( .D(n2943), .CK(n993), .QN(n672) );
  DFF_X1 \reg_22/q_reg[0]  ( .D(n2942), .CK(n993), .QN(n673) );
  DFF_X1 \reg_22/q_reg[1]  ( .D(n2941), .CK(n993), .QN(n674) );
  DFF_X1 \reg_22/q_reg[2]  ( .D(n2940), .CK(n993), .QN(n675) );
  DFF_X1 \reg_22/q_reg[3]  ( .D(n2939), .CK(n993), .QN(n676) );
  DFF_X1 \reg_22/q_reg[4]  ( .D(n2938), .CK(n993), .QN(n677) );
  DFF_X1 \reg_22/q_reg[5]  ( .D(n2937), .CK(n993), .QN(n678) );
  DFF_X1 \reg_22/q_reg[6]  ( .D(n2936), .CK(n993), .QN(n679) );
  DFF_X1 \reg_22/q_reg[7]  ( .D(n2935), .CK(n993), .QN(n680) );
  DFF_X1 \reg_22/q_reg[8]  ( .D(n2934), .CK(n993), .QN(n681) );
  DFF_X1 \reg_22/q_reg[9]  ( .D(n2933), .CK(n993), .QN(n682) );
  DFF_X1 \reg_22/q_reg[10]  ( .D(n2932), .CK(n993), .QN(n683) );
  DFF_X1 \reg_22/q_reg[11]  ( .D(n2931), .CK(n993), .QN(n684) );
  DFF_X1 \reg_22/q_reg[12]  ( .D(n2930), .CK(n993), .QN(n685) );
  DFF_X1 \reg_22/q_reg[13]  ( .D(n2929), .CK(n993), .QN(n686) );
  DFF_X1 \reg_22/q_reg[14]  ( .D(n2928), .CK(n993), .QN(n687) );
  DFF_X1 \reg_22/q_reg[15]  ( .D(n2927), .CK(n993), .QN(n688) );
  DFF_X1 \reg_22/q_reg[16]  ( .D(n2926), .CK(n993), .QN(n689) );
  DFF_X1 \reg_22/q_reg[17]  ( .D(n2925), .CK(n993), .QN(n690) );
  DFF_X1 \reg_22/q_reg[18]  ( .D(n2924), .CK(n993), .QN(n691) );
  DFF_X1 \reg_22/q_reg[19]  ( .D(n2923), .CK(n993), .QN(n692) );
  DFF_X1 \reg_22/q_reg[20]  ( .D(n2922), .CK(n993), .QN(n693) );
  DFF_X1 \reg_22/q_reg[21]  ( .D(n2921), .CK(n993), .QN(n694) );
  DFF_X1 \reg_22/q_reg[22]  ( .D(n2920), .CK(n993), .QN(n695) );
  DFF_X1 \reg_22/q_reg[23]  ( .D(n2919), .CK(n993), .QN(n696) );
  DFF_X1 \reg_22/q_reg[24]  ( .D(n2918), .CK(n993), .QN(n697) );
  DFF_X1 \reg_22/q_reg[25]  ( .D(n2917), .CK(n993), .QN(n698) );
  DFF_X1 \reg_22/q_reg[26]  ( .D(n2916), .CK(n993), .QN(n699) );
  DFF_X1 \reg_22/q_reg[27]  ( .D(n2915), .CK(n993), .QN(n700) );
  DFF_X1 \reg_22/q_reg[28]  ( .D(n2914), .CK(n993), .QN(n701) );
  DFF_X1 \reg_22/q_reg[29]  ( .D(n2913), .CK(n993), .QN(n702) );
  DFF_X1 \reg_22/q_reg[30]  ( .D(n2912), .CK(n993), .QN(n703) );
  DFF_X1 \reg_22/q_reg[31]  ( .D(n2911), .CK(n993), .QN(n704) );
  DFF_X1 \reg_23/q_reg[0]  ( .D(n2910), .CK(n993), .QN(n705) );
  DFF_X1 \reg_23/q_reg[1]  ( .D(n2909), .CK(n993), .QN(n706) );
  DFF_X1 \reg_23/q_reg[2]  ( .D(n2908), .CK(n993), .QN(n707) );
  DFF_X1 \reg_23/q_reg[3]  ( .D(n2907), .CK(n993), .QN(n708) );
  DFF_X1 \reg_23/q_reg[4]  ( .D(n2906), .CK(n993), .QN(n709) );
  DFF_X1 \reg_23/q_reg[5]  ( .D(n2905), .CK(n993), .QN(n710) );
  DFF_X1 \reg_23/q_reg[6]  ( .D(n2904), .CK(n993), .QN(n711) );
  DFF_X1 \reg_23/q_reg[7]  ( .D(n2903), .CK(n993), .QN(n712) );
  DFF_X1 \reg_23/q_reg[8]  ( .D(n2902), .CK(n993), .QN(n713) );
  DFF_X1 \reg_23/q_reg[9]  ( .D(n2901), .CK(n993), .QN(n714) );
  DFF_X1 \reg_23/q_reg[10]  ( .D(n2900), .CK(n993), .QN(n715) );
  DFF_X1 \reg_23/q_reg[11]  ( .D(n2899), .CK(n993), .QN(n716) );
  DFF_X1 \reg_23/q_reg[12]  ( .D(n2898), .CK(n993), .QN(n717) );
  DFF_X1 \reg_23/q_reg[13]  ( .D(n2897), .CK(n993), .QN(n718) );
  DFF_X1 \reg_23/q_reg[14]  ( .D(n2896), .CK(n993), .QN(n719) );
  DFF_X1 \reg_23/q_reg[15]  ( .D(n2895), .CK(n993), .QN(n720) );
  DFF_X1 \reg_23/q_reg[16]  ( .D(n2894), .CK(n993), .QN(n721) );
  DFF_X1 \reg_23/q_reg[17]  ( .D(n2893), .CK(n993), .QN(n722) );
  DFF_X1 \reg_23/q_reg[18]  ( .D(n2892), .CK(n993), .QN(n723) );
  DFF_X1 \reg_23/q_reg[19]  ( .D(n2891), .CK(n993), .QN(n724) );
  DFF_X1 \reg_23/q_reg[20]  ( .D(n2890), .CK(n993), .QN(n725) );
  DFF_X1 \reg_23/q_reg[21]  ( .D(n2889), .CK(n993), .QN(n726) );
  DFF_X1 \reg_23/q_reg[22]  ( .D(n2888), .CK(n993), .QN(n727) );
  DFF_X1 \reg_23/q_reg[23]  ( .D(n2887), .CK(n993), .QN(n728) );
  DFF_X1 \reg_23/q_reg[24]  ( .D(n2886), .CK(n993), .QN(n729) );
  DFF_X1 \reg_23/q_reg[25]  ( .D(n2885), .CK(n993), .QN(n730) );
  DFF_X1 \reg_23/q_reg[26]  ( .D(n2884), .CK(n993), .QN(n731) );
  DFF_X1 \reg_23/q_reg[27]  ( .D(n2883), .CK(n993), .QN(n732) );
  DFF_X1 \reg_23/q_reg[28]  ( .D(n2882), .CK(n993), .QN(n733) );
  DFF_X1 \reg_23/q_reg[29]  ( .D(n2881), .CK(n993), .QN(n734) );
  DFF_X1 \reg_23/q_reg[30]  ( .D(n2880), .CK(n993), .QN(n735) );
  DFF_X1 \reg_23/q_reg[31]  ( .D(n2879), .CK(n993), .QN(n736) );
  DFF_X1 \reg_24/q_reg[0]  ( .D(n2878), .CK(n993), .QN(n737) );
  DFF_X1 \reg_24/q_reg[1]  ( .D(n2877), .CK(n993), .QN(n738) );
  DFF_X1 \reg_24/q_reg[2]  ( .D(n2876), .CK(n993), .QN(n739) );
  DFF_X1 \reg_24/q_reg[3]  ( .D(n2875), .CK(n993), .QN(n740) );
  DFF_X1 \reg_24/q_reg[4]  ( .D(n2874), .CK(n993), .QN(n741) );
  DFF_X1 \reg_24/q_reg[5]  ( .D(n2873), .CK(n993), .QN(n742) );
  DFF_X1 \reg_24/q_reg[6]  ( .D(n2872), .CK(n993), .QN(n743) );
  DFF_X1 \reg_24/q_reg[7]  ( .D(n2871), .CK(n993), .QN(n744) );
  DFF_X1 \reg_24/q_reg[8]  ( .D(n2870), .CK(n993), .QN(n745) );
  DFF_X1 \reg_24/q_reg[9]  ( .D(n2869), .CK(n993), .QN(n746) );
  DFF_X1 \reg_24/q_reg[10]  ( .D(n2868), .CK(n993), .QN(n747) );
  DFF_X1 \reg_24/q_reg[11]  ( .D(n2867), .CK(n993), .QN(n748) );
  DFF_X1 \reg_24/q_reg[12]  ( .D(n2866), .CK(n993), .QN(n749) );
  DFF_X1 \reg_24/q_reg[13]  ( .D(n2865), .CK(n993), .QN(n750) );
  DFF_X1 \reg_24/q_reg[14]  ( .D(n2864), .CK(n993), .QN(n751) );
  DFF_X1 \reg_24/q_reg[15]  ( .D(n2863), .CK(n993), .QN(n752) );
  DFF_X1 \reg_24/q_reg[16]  ( .D(n2862), .CK(n993), .QN(n753) );
  DFF_X1 \reg_24/q_reg[17]  ( .D(n2861), .CK(n993), .QN(n754) );
  DFF_X1 \reg_24/q_reg[18]  ( .D(n2860), .CK(n993), .QN(n755) );
  DFF_X1 \reg_24/q_reg[19]  ( .D(n2859), .CK(n993), .QN(n756) );
  DFF_X1 \reg_24/q_reg[20]  ( .D(n2858), .CK(n993), .QN(n757) );
  DFF_X1 \reg_24/q_reg[21]  ( .D(n2857), .CK(n993), .QN(n758) );
  DFF_X1 \reg_24/q_reg[22]  ( .D(n2856), .CK(n993), .QN(n759) );
  DFF_X1 \reg_24/q_reg[23]  ( .D(n2855), .CK(n993), .QN(n760) );
  DFF_X1 \reg_24/q_reg[24]  ( .D(n2854), .CK(n993), .QN(n761) );
  DFF_X1 \reg_24/q_reg[25]  ( .D(n2853), .CK(n993), .QN(n762) );
  DFF_X1 \reg_24/q_reg[26]  ( .D(n2852), .CK(n993), .QN(n763) );
  DFF_X1 \reg_24/q_reg[27]  ( .D(n2851), .CK(n993), .QN(n764) );
  DFF_X1 \reg_24/q_reg[28]  ( .D(n2850), .CK(n993), .QN(n765) );
  DFF_X1 \reg_24/q_reg[29]  ( .D(n2849), .CK(n993), .QN(n766) );
  DFF_X1 \reg_24/q_reg[30]  ( .D(n2848), .CK(n993), .QN(n767) );
  DFF_X1 \reg_24/q_reg[31]  ( .D(n2847), .CK(n993), .QN(n768) );
  DFF_X1 \reg_25/q_reg[0]  ( .D(n2846), .CK(n993), .QN(n769) );
  DFF_X1 \reg_25/q_reg[1]  ( .D(n2845), .CK(n993), .QN(n770) );
  DFF_X1 \reg_25/q_reg[2]  ( .D(n2844), .CK(n993), .QN(n771) );
  DFF_X1 \reg_25/q_reg[3]  ( .D(n2843), .CK(n993), .QN(n772) );
  DFF_X1 \reg_25/q_reg[4]  ( .D(n2842), .CK(n993), .QN(n773) );
  DFF_X1 \reg_25/q_reg[5]  ( .D(n2841), .CK(n993), .QN(n774) );
  DFF_X1 \reg_25/q_reg[6]  ( .D(n2840), .CK(n993), .QN(n775) );
  DFF_X1 \reg_25/q_reg[7]  ( .D(n2839), .CK(n993), .QN(n776) );
  DFF_X1 \reg_25/q_reg[8]  ( .D(n2838), .CK(n993), .QN(n777) );
  DFF_X1 \reg_25/q_reg[9]  ( .D(n2837), .CK(n993), .QN(n778) );
  DFF_X1 \reg_25/q_reg[10]  ( .D(n2836), .CK(n993), .QN(n779) );
  DFF_X1 \reg_25/q_reg[11]  ( .D(n2835), .CK(n993), .QN(n780) );
  DFF_X1 \reg_25/q_reg[12]  ( .D(n2834), .CK(n993), .QN(n781) );
  DFF_X1 \reg_25/q_reg[13]  ( .D(n2833), .CK(n993), .QN(n782) );
  DFF_X1 \reg_25/q_reg[14]  ( .D(n2832), .CK(n993), .QN(n783) );
  DFF_X1 \reg_25/q_reg[15]  ( .D(n2831), .CK(n993), .QN(n784) );
  DFF_X1 \reg_25/q_reg[16]  ( .D(n2830), .CK(n993), .QN(n785) );
  DFF_X1 \reg_25/q_reg[17]  ( .D(n2829), .CK(n993), .QN(n786) );
  DFF_X1 \reg_25/q_reg[18]  ( .D(n2828), .CK(n993), .QN(n787) );
  DFF_X1 \reg_25/q_reg[19]  ( .D(n2827), .CK(n993), .QN(n788) );
  DFF_X1 \reg_25/q_reg[20]  ( .D(n2826), .CK(n993), .QN(n789) );
  DFF_X1 \reg_25/q_reg[21]  ( .D(n2825), .CK(n993), .QN(n790) );
  DFF_X1 \reg_25/q_reg[22]  ( .D(n2824), .CK(n993), .QN(n791) );
  DFF_X1 \reg_25/q_reg[23]  ( .D(n2823), .CK(n993), .QN(n792) );
  DFF_X1 \reg_25/q_reg[24]  ( .D(n2822), .CK(n993), .QN(n793) );
  DFF_X1 \reg_25/q_reg[25]  ( .D(n2821), .CK(n993), .QN(n794) );
  DFF_X1 \reg_25/q_reg[26]  ( .D(n2820), .CK(n993), .QN(n795) );
  DFF_X1 \reg_25/q_reg[27]  ( .D(n2819), .CK(n993), .QN(n796) );
  DFF_X1 \reg_25/q_reg[28]  ( .D(n2818), .CK(n993), .QN(n797) );
  DFF_X1 \reg_25/q_reg[29]  ( .D(n2817), .CK(n993), .QN(n798) );
  DFF_X1 \reg_25/q_reg[30]  ( .D(n2816), .CK(n993), .QN(n799) );
  DFF_X1 \reg_25/q_reg[31]  ( .D(n2815), .CK(n993), .QN(n800) );
  DFF_X1 \reg_26/q_reg[0]  ( .D(n2814), .CK(n993), .QN(n801) );
  DFF_X1 \reg_26/q_reg[1]  ( .D(n2813), .CK(n993), .QN(n802) );
  DFF_X1 \reg_26/q_reg[2]  ( .D(n2812), .CK(n993), .QN(n803) );
  DFF_X1 \reg_26/q_reg[3]  ( .D(n2811), .CK(n993), .QN(n804) );
  DFF_X1 \reg_26/q_reg[4]  ( .D(n2810), .CK(n993), .QN(n805) );
  DFF_X1 \reg_26/q_reg[5]  ( .D(n2809), .CK(n993), .QN(n806) );
  DFF_X1 \reg_26/q_reg[6]  ( .D(n2808), .CK(n993), .QN(n807) );
  DFF_X1 \reg_26/q_reg[7]  ( .D(n2807), .CK(n993), .QN(n808) );
  DFF_X1 \reg_26/q_reg[8]  ( .D(n2806), .CK(n993), .QN(n809) );
  DFF_X1 \reg_26/q_reg[9]  ( .D(n2805), .CK(n993), .QN(n810) );
  DFF_X1 \reg_26/q_reg[10]  ( .D(n2804), .CK(n993), .QN(n811) );
  DFF_X1 \reg_26/q_reg[11]  ( .D(n2803), .CK(n993), .QN(n812) );
  DFF_X1 \reg_26/q_reg[12]  ( .D(n2802), .CK(n993), .QN(n813) );
  DFF_X1 \reg_26/q_reg[13]  ( .D(n2801), .CK(n993), .QN(n814) );
  DFF_X1 \reg_26/q_reg[14]  ( .D(n2800), .CK(n993), .QN(n815) );
  DFF_X1 \reg_26/q_reg[15]  ( .D(n2799), .CK(n993), .QN(n816) );
  DFF_X1 \reg_26/q_reg[16]  ( .D(n2798), .CK(n993), .QN(n817) );
  DFF_X1 \reg_26/q_reg[17]  ( .D(n2797), .CK(n993), .QN(n818) );
  DFF_X1 \reg_26/q_reg[18]  ( .D(n2796), .CK(n993), .QN(n819) );
  DFF_X1 \reg_26/q_reg[19]  ( .D(n2795), .CK(n993), .QN(n820) );
  DFF_X1 \reg_26/q_reg[20]  ( .D(n2794), .CK(n993), .QN(n821) );
  DFF_X1 \reg_26/q_reg[21]  ( .D(n2793), .CK(n993), .QN(n822) );
  DFF_X1 \reg_26/q_reg[22]  ( .D(n2792), .CK(n993), .QN(n823) );
  DFF_X1 \reg_26/q_reg[23]  ( .D(n2791), .CK(n993), .QN(n824) );
  DFF_X1 \reg_26/q_reg[24]  ( .D(n2790), .CK(n993), .QN(n825) );
  DFF_X1 \reg_26/q_reg[25]  ( .D(n2789), .CK(n993), .QN(n826) );
  DFF_X1 \reg_26/q_reg[26]  ( .D(n2788), .CK(n993), .QN(n827) );
  DFF_X1 \reg_26/q_reg[27]  ( .D(n2787), .CK(n993), .QN(n828) );
  DFF_X1 \reg_26/q_reg[28]  ( .D(n2786), .CK(n993), .QN(n829) );
  DFF_X1 \reg_26/q_reg[29]  ( .D(n2785), .CK(n993), .QN(n830) );
  DFF_X1 \reg_26/q_reg[30]  ( .D(n2784), .CK(n993), .QN(n831) );
  DFF_X1 \reg_26/q_reg[31]  ( .D(n2783), .CK(n993), .QN(n832) );
  DFF_X1 \reg_27/q_reg[0]  ( .D(n2782), .CK(n993), .QN(n833) );
  DFF_X1 \reg_27/q_reg[1]  ( .D(n2781), .CK(n993), .QN(n834) );
  DFF_X1 \reg_27/q_reg[2]  ( .D(n2780), .CK(n993), .QN(n835) );
  DFF_X1 \reg_27/q_reg[3]  ( .D(n2779), .CK(n993), .QN(n836) );
  DFF_X1 \reg_27/q_reg[4]  ( .D(n2778), .CK(n993), .QN(n837) );
  DFF_X1 \reg_27/q_reg[5]  ( .D(n2777), .CK(n993), .QN(n838) );
  DFF_X1 \reg_27/q_reg[6]  ( .D(n2776), .CK(n993), .QN(n839) );
  DFF_X1 \reg_27/q_reg[7]  ( .D(n2775), .CK(n993), .QN(n840) );
  DFF_X1 \reg_27/q_reg[8]  ( .D(n2774), .CK(n993), .QN(n841) );
  DFF_X1 \reg_27/q_reg[9]  ( .D(n2773), .CK(n993), .QN(n842) );
  DFF_X1 \reg_27/q_reg[10]  ( .D(n2772), .CK(n993), .QN(n843) );
  DFF_X1 \reg_27/q_reg[11]  ( .D(n2771), .CK(n993), .QN(n844) );
  DFF_X1 \reg_27/q_reg[12]  ( .D(n2770), .CK(n993), .QN(n845) );
  DFF_X1 \reg_27/q_reg[13]  ( .D(n2769), .CK(n993), .QN(n846) );
  DFF_X1 \reg_27/q_reg[14]  ( .D(n2768), .CK(n993), .QN(n847) );
  DFF_X1 \reg_27/q_reg[15]  ( .D(n2767), .CK(n993), .QN(n848) );
  DFF_X1 \reg_27/q_reg[16]  ( .D(n2766), .CK(n993), .QN(n849) );
  DFF_X1 \reg_27/q_reg[17]  ( .D(n2765), .CK(n993), .QN(n850) );
  DFF_X1 \reg_27/q_reg[18]  ( .D(n2764), .CK(n993), .QN(n851) );
  DFF_X1 \reg_27/q_reg[19]  ( .D(n2763), .CK(n993), .QN(n852) );
  DFF_X1 \reg_27/q_reg[20]  ( .D(n2762), .CK(n993), .QN(n853) );
  DFF_X1 \reg_27/q_reg[21]  ( .D(n2761), .CK(n993), .QN(n854) );
  DFF_X1 \reg_27/q_reg[22]  ( .D(n2760), .CK(n993), .QN(n855) );
  DFF_X1 \reg_27/q_reg[23]  ( .D(n2759), .CK(n993), .QN(n856) );
  DFF_X1 \reg_27/q_reg[24]  ( .D(n2758), .CK(n993), .QN(n857) );
  DFF_X1 \reg_27/q_reg[25]  ( .D(n2757), .CK(n993), .QN(n858) );
  DFF_X1 \reg_27/q_reg[26]  ( .D(n2756), .CK(n993), .QN(n859) );
  DFF_X1 \reg_27/q_reg[27]  ( .D(n2755), .CK(n993), .QN(n860) );
  DFF_X1 \reg_27/q_reg[28]  ( .D(n2754), .CK(n993), .QN(n861) );
  DFF_X1 \reg_27/q_reg[29]  ( .D(n2753), .CK(n993), .QN(n862) );
  DFF_X1 \reg_27/q_reg[30]  ( .D(n2752), .CK(n993), .QN(n863) );
  DFF_X1 \reg_27/q_reg[31]  ( .D(n2751), .CK(n993), .QN(n864) );
  DFF_X1 \reg_28/q_reg[0]  ( .D(n2750), .CK(n993), .QN(n865) );
  DFF_X1 \reg_28/q_reg[1]  ( .D(n2749), .CK(n993), .QN(n866) );
  DFF_X1 \reg_28/q_reg[2]  ( .D(n2748), .CK(n993), .QN(n867) );
  DFF_X1 \reg_28/q_reg[3]  ( .D(n2747), .CK(n993), .QN(n868) );
  DFF_X1 \reg_28/q_reg[4]  ( .D(n2746), .CK(n993), .QN(n869) );
  DFF_X1 \reg_28/q_reg[5]  ( .D(n2745), .CK(n993), .QN(n870) );
  DFF_X1 \reg_28/q_reg[6]  ( .D(n2744), .CK(n993), .QN(n871) );
  DFF_X1 \reg_28/q_reg[7]  ( .D(n2743), .CK(n993), .QN(n872) );
  DFF_X1 \reg_28/q_reg[8]  ( .D(n2742), .CK(n993), .QN(n873) );
  DFF_X1 \reg_28/q_reg[9]  ( .D(n2741), .CK(n993), .QN(n874) );
  DFF_X1 \reg_28/q_reg[10]  ( .D(n2740), .CK(n993), .QN(n875) );
  DFF_X1 \reg_28/q_reg[11]  ( .D(n2739), .CK(n993), .QN(n876) );
  DFF_X1 \reg_28/q_reg[12]  ( .D(n2738), .CK(n993), .QN(n877) );
  DFF_X1 \reg_28/q_reg[13]  ( .D(n2737), .CK(n993), .QN(n878) );
  DFF_X1 \reg_28/q_reg[14]  ( .D(n2736), .CK(n993), .QN(n879) );
  DFF_X1 \reg_28/q_reg[15]  ( .D(n2735), .CK(n993), .QN(n880) );
  DFF_X1 \reg_28/q_reg[16]  ( .D(n2734), .CK(n993), .QN(n881) );
  DFF_X1 \reg_28/q_reg[17]  ( .D(n2733), .CK(n993), .QN(n882) );
  DFF_X1 \reg_28/q_reg[18]  ( .D(n2732), .CK(n993), .QN(n883) );
  DFF_X1 \reg_28/q_reg[19]  ( .D(n2731), .CK(n993), .QN(n884) );
  DFF_X1 \reg_28/q_reg[20]  ( .D(n2730), .CK(n993), .QN(n885) );
  DFF_X1 \reg_28/q_reg[21]  ( .D(n2729), .CK(n993), .QN(n886) );
  DFF_X1 \reg_28/q_reg[22]  ( .D(n2728), .CK(n993), .QN(n887) );
  DFF_X1 \reg_28/q_reg[23]  ( .D(n2727), .CK(n993), .QN(n888) );
  DFF_X1 \reg_28/q_reg[24]  ( .D(n2726), .CK(n993), .QN(n889) );
  DFF_X1 \reg_28/q_reg[25]  ( .D(n2725), .CK(n993), .QN(n890) );
  DFF_X1 \reg_28/q_reg[26]  ( .D(n2724), .CK(n993), .QN(n891) );
  DFF_X1 \reg_28/q_reg[27]  ( .D(n2723), .CK(n993), .QN(n892) );
  DFF_X1 \reg_28/q_reg[28]  ( .D(n2722), .CK(n993), .QN(n893) );
  DFF_X1 \reg_28/q_reg[29]  ( .D(n2721), .CK(n993), .QN(n894) );
  DFF_X1 \reg_28/q_reg[30]  ( .D(n2720), .CK(n993), .QN(n895) );
  DFF_X1 \reg_28/q_reg[31]  ( .D(n2719), .CK(n993), .QN(n896) );
  DFF_X1 \reg_29/q_reg[0]  ( .D(n2718), .CK(n993), .QN(n897) );
  DFF_X1 \reg_29/q_reg[1]  ( .D(n2717), .CK(n993), .QN(n898) );
  DFF_X1 \reg_29/q_reg[2]  ( .D(n2716), .CK(n993), .QN(n899) );
  DFF_X1 \reg_29/q_reg[3]  ( .D(n2715), .CK(n993), .QN(n900) );
  DFF_X1 \reg_29/q_reg[4]  ( .D(n2714), .CK(n993), .QN(n901) );
  DFF_X1 \reg_29/q_reg[5]  ( .D(n2713), .CK(n993), .QN(n902) );
  DFF_X1 \reg_29/q_reg[6]  ( .D(n2712), .CK(n993), .QN(n903) );
  DFF_X1 \reg_29/q_reg[7]  ( .D(n2711), .CK(n993), .QN(n904) );
  DFF_X1 \reg_29/q_reg[8]  ( .D(n2710), .CK(n993), .QN(n905) );
  DFF_X1 \reg_29/q_reg[9]  ( .D(n2709), .CK(n993), .QN(n906) );
  DFF_X1 \reg_29/q_reg[10]  ( .D(n2708), .CK(n993), .QN(n907) );
  DFF_X1 \reg_29/q_reg[11]  ( .D(n2707), .CK(n993), .QN(n908) );
  DFF_X1 \reg_29/q_reg[12]  ( .D(n2706), .CK(n993), .QN(n909) );
  DFF_X1 \reg_29/q_reg[13]  ( .D(n2705), .CK(n993), .QN(n910) );
  DFF_X1 \reg_29/q_reg[14]  ( .D(n2704), .CK(n993), .QN(n911) );
  DFF_X1 \reg_29/q_reg[15]  ( .D(n2703), .CK(n993), .QN(n912) );
  DFF_X1 \reg_29/q_reg[16]  ( .D(n2702), .CK(n993), .QN(n913) );
  DFF_X1 \reg_29/q_reg[17]  ( .D(n2701), .CK(n993), .QN(n914) );
  DFF_X1 \reg_29/q_reg[18]  ( .D(n2700), .CK(n993), .QN(n915) );
  DFF_X1 \reg_29/q_reg[19]  ( .D(n2699), .CK(n993), .QN(n916) );
  DFF_X1 \reg_29/q_reg[20]  ( .D(n2698), .CK(n993), .QN(n917) );
  DFF_X1 \reg_29/q_reg[21]  ( .D(n2697), .CK(n993), .QN(n918) );
  DFF_X1 \reg_29/q_reg[22]  ( .D(n2696), .CK(n993), .QN(n919) );
  DFF_X1 \reg_29/q_reg[23]  ( .D(n2695), .CK(n993), .QN(n920) );
  DFF_X1 \reg_29/q_reg[24]  ( .D(n2694), .CK(n993), .QN(n921) );
  DFF_X1 \reg_29/q_reg[25]  ( .D(n2693), .CK(n993), .QN(n922) );
  DFF_X1 \reg_29/q_reg[26]  ( .D(n2692), .CK(n993), .QN(n923) );
  DFF_X1 \reg_29/q_reg[27]  ( .D(n2691), .CK(n993), .QN(n924) );
  DFF_X1 \reg_29/q_reg[28]  ( .D(n2690), .CK(n993), .QN(n925) );
  DFF_X1 \reg_29/q_reg[29]  ( .D(n2689), .CK(n993), .QN(n926) );
  DFF_X1 \reg_29/q_reg[30]  ( .D(n2688), .CK(n993), .QN(n927) );
  DFF_X1 \reg_29/q_reg[31]  ( .D(n2687), .CK(n993), .QN(n928) );
  DFF_X1 \reg_30/q_reg[0]  ( .D(n2686), .CK(n993), .QN(n929) );
  DFF_X1 \reg_30/q_reg[1]  ( .D(n2685), .CK(n993), .QN(n930) );
  DFF_X1 \reg_30/q_reg[2]  ( .D(n2684), .CK(n993), .QN(n931) );
  DFF_X1 \reg_30/q_reg[3]  ( .D(n2683), .CK(n993), .QN(n932) );
  DFF_X1 \reg_30/q_reg[4]  ( .D(n2682), .CK(n993), .QN(n933) );
  DFF_X1 \reg_30/q_reg[5]  ( .D(n2681), .CK(n993), .QN(n934) );
  DFF_X1 \reg_30/q_reg[6]  ( .D(n2680), .CK(n993), .QN(n935) );
  DFF_X1 \reg_30/q_reg[7]  ( .D(n2679), .CK(n993), .QN(n936) );
  DFF_X1 \reg_30/q_reg[8]  ( .D(n2678), .CK(n993), .QN(n937) );
  DFF_X1 \reg_30/q_reg[9]  ( .D(n2677), .CK(n993), .QN(n938) );
  DFF_X1 \reg_30/q_reg[10]  ( .D(n2676), .CK(n993), .QN(n939) );
  DFF_X1 \reg_30/q_reg[11]  ( .D(n2675), .CK(n993), .QN(n940) );
  DFF_X1 \reg_30/q_reg[12]  ( .D(n2674), .CK(n993), .QN(n941) );
  DFF_X1 \reg_30/q_reg[13]  ( .D(n2673), .CK(n993), .QN(n942) );
  DFF_X1 \reg_30/q_reg[14]  ( .D(n2672), .CK(n993), .QN(n943) );
  DFF_X1 \reg_30/q_reg[15]  ( .D(n2671), .CK(n993), .QN(n944) );
  DFF_X1 \reg_30/q_reg[16]  ( .D(n2670), .CK(n993), .QN(n945) );
  DFF_X1 \reg_30/q_reg[17]  ( .D(n2669), .CK(n993), .QN(n946) );
  DFF_X1 \reg_30/q_reg[18]  ( .D(n2668), .CK(n993), .QN(n947) );
  DFF_X1 \reg_30/q_reg[19]  ( .D(n2667), .CK(n993), .QN(n948) );
  DFF_X1 \reg_30/q_reg[20]  ( .D(n2666), .CK(n993), .QN(n949) );
  DFF_X1 \reg_30/q_reg[21]  ( .D(n2665), .CK(n993), .QN(n950) );
  DFF_X1 \reg_30/q_reg[22]  ( .D(n2664), .CK(n993), .QN(n951) );
  DFF_X1 \reg_30/q_reg[23]  ( .D(n2663), .CK(n993), .QN(n952) );
  DFF_X1 \reg_30/q_reg[24]  ( .D(n2662), .CK(n993), .QN(n953) );
  DFF_X1 \reg_30/q_reg[25]  ( .D(n2661), .CK(n993), .QN(n954) );
  DFF_X1 \reg_30/q_reg[26]  ( .D(n2660), .CK(n993), .QN(n955) );
  DFF_X1 \reg_30/q_reg[27]  ( .D(n2659), .CK(n993), .QN(n956) );
  DFF_X1 \reg_30/q_reg[28]  ( .D(n2658), .CK(n993), .QN(n957) );
  DFF_X1 \reg_30/q_reg[29]  ( .D(n2657), .CK(n993), .QN(n958) );
  DFF_X1 \reg_30/q_reg[30]  ( .D(n2656), .CK(n993), .QN(n959) );
  DFF_X1 \reg_30/q_reg[31]  ( .D(n2655), .CK(n993), .QN(n960) );
  DFF_X1 \reg_31/q_reg[0]  ( .D(n2654), .CK(n993), .QN(n961) );
  DFF_X1 \reg_31/q_reg[1]  ( .D(n2653), .CK(n993), .QN(n962) );
  DFF_X1 \reg_31/q_reg[2]  ( .D(n2652), .CK(n993), .QN(n963) );
  DFF_X1 \reg_31/q_reg[3]  ( .D(n2651), .CK(n993), .QN(n964) );
  DFF_X1 \reg_31/q_reg[4]  ( .D(n2650), .CK(n993), .QN(n965) );
  DFF_X1 \reg_31/q_reg[5]  ( .D(n2649), .CK(n993), .QN(n966) );
  DFF_X1 \reg_31/q_reg[6]  ( .D(n2648), .CK(n993), .QN(n967) );
  DFF_X1 \reg_31/q_reg[7]  ( .D(n2647), .CK(n993), .QN(n968) );
  DFF_X1 \reg_31/q_reg[8]  ( .D(n2646), .CK(n993), .QN(n969) );
  DFF_X1 \reg_31/q_reg[9]  ( .D(n2645), .CK(n993), .QN(n970) );
  DFF_X1 \reg_31/q_reg[10]  ( .D(n2644), .CK(n993), .QN(n971) );
  DFF_X1 \reg_31/q_reg[11]  ( .D(n2643), .CK(n993), .QN(n972) );
  DFF_X1 \reg_31/q_reg[12]  ( .D(n2642), .CK(n993), .QN(n973) );
  DFF_X1 \reg_31/q_reg[13]  ( .D(n2641), .CK(n993), .QN(n974) );
  DFF_X1 \reg_31/q_reg[14]  ( .D(n2640), .CK(n993), .QN(n975) );
  DFF_X1 \reg_31/q_reg[15]  ( .D(n2639), .CK(n993), .QN(n976) );
  DFF_X1 \reg_31/q_reg[16]  ( .D(n2638), .CK(n993), .QN(n977) );
  DFF_X1 \reg_31/q_reg[17]  ( .D(n2637), .CK(n993), .QN(n978) );
  DFF_X1 \reg_31/q_reg[18]  ( .D(n2636), .CK(n993), .QN(n979) );
  DFF_X1 \reg_31/q_reg[19]  ( .D(n2635), .CK(n993), .QN(n980) );
  DFF_X1 \reg_31/q_reg[20]  ( .D(n2634), .CK(n993), .QN(n981) );
  DFF_X1 \reg_31/q_reg[21]  ( .D(n2633), .CK(n993), .QN(n982) );
  DFF_X1 \reg_31/q_reg[22]  ( .D(n2632), .CK(n993), .QN(n983) );
  DFF_X1 \reg_31/q_reg[23]  ( .D(n2631), .CK(n993), .QN(n984) );
  DFF_X1 \reg_31/q_reg[24]  ( .D(n2630), .CK(n993), .QN(n985) );
  DFF_X1 \reg_31/q_reg[25]  ( .D(n2629), .CK(n993), .QN(n986) );
  DFF_X1 \reg_31/q_reg[26]  ( .D(n2628), .CK(n993), .QN(n987) );
  DFF_X1 \reg_31/q_reg[27]  ( .D(n2627), .CK(n993), .QN(n988) );
  DFF_X1 \reg_31/q_reg[28]  ( .D(n2626), .CK(n993), .QN(n989) );
  DFF_X1 \reg_31/q_reg[29]  ( .D(n2625), .CK(n993), .QN(n990) );
  DFF_X1 \reg_31/q_reg[30]  ( .D(n2624), .CK(n993), .QN(n991) );
  DFF_X1 \reg_31/q_reg[31]  ( .D(n2623), .CK(n993), .QN(n992) );
  DFF_X1 \lo/q_reg[0]  ( .D(n2547), .CK(n993), .QN(lo_out[0]) );
  DFF_X1 \lo/q_reg[1]  ( .D(n2546), .CK(n993), .QN(lo_out[1]) );
  DFF_X1 \lo/q_reg[2]  ( .D(n2545), .CK(n993), .QN(lo_out[2]) );
  DFF_X1 \lo/q_reg[3]  ( .D(n2544), .CK(n993), .QN(lo_out[3]) );
  DFF_X1 \lo/q_reg[4]  ( .D(n2543), .CK(n993), .QN(lo_out[4]) );
  DFF_X1 \lo/q_reg[5]  ( .D(n2542), .CK(n993), .QN(lo_out[5]) );
  DFF_X1 \lo/q_reg[6]  ( .D(n2541), .CK(n993), .QN(lo_out[6]) );
  DFF_X1 \lo/q_reg[7]  ( .D(n2540), .CK(n993), .QN(lo_out[7]) );
  DFF_X1 \lo/q_reg[8]  ( .D(n2539), .CK(n993), .QN(lo_out[8]) );
  DFF_X1 \lo/q_reg[9]  ( .D(n2538), .CK(n993), .QN(lo_out[9]) );
  DFF_X1 \lo/q_reg[10]  ( .D(n2537), .CK(n993), .QN(lo_out[10]) );
  DFF_X1 \lo/q_reg[11]  ( .D(n2536), .CK(n993), .QN(lo_out[11]) );
  DFF_X1 \lo/q_reg[12]  ( .D(n2535), .CK(n993), .QN(lo_out[12]) );
  DFF_X1 \lo/q_reg[13]  ( .D(n2534), .CK(n993), .QN(lo_out[13]) );
  DFF_X1 \lo/q_reg[14]  ( .D(n2533), .CK(n993), .QN(lo_out[14]) );
  DFF_X1 \lo/q_reg[15]  ( .D(n2532), .CK(n993), .QN(lo_out[15]) );
  DFF_X1 \lo/q_reg[16]  ( .D(n2531), .CK(n993), .QN(lo_out[16]) );
  DFF_X1 \lo/q_reg[17]  ( .D(n2530), .CK(n993), .QN(lo_out[17]) );
  DFF_X1 \lo/q_reg[18]  ( .D(n2529), .CK(n993), .QN(lo_out[18]) );
  DFF_X1 \lo/q_reg[19]  ( .D(n2528), .CK(n993), .QN(lo_out[19]) );
  DFF_X1 \lo/q_reg[20]  ( .D(n2527), .CK(n993), .QN(lo_out[20]) );
  DFF_X1 \lo/q_reg[21]  ( .D(n2526), .CK(n993), .QN(lo_out[21]) );
  DFF_X1 \lo/q_reg[22]  ( .D(n2525), .CK(n993), .QN(lo_out[22]) );
  DFF_X1 \lo/q_reg[23]  ( .D(n2524), .CK(n993), .QN(lo_out[23]) );
  DFF_X1 \lo/q_reg[24]  ( .D(n2523), .CK(n993), .QN(lo_out[24]) );
  DFF_X1 \lo/q_reg[25]  ( .D(n2522), .CK(n993), .QN(lo_out[25]) );
  DFF_X1 \lo/q_reg[26]  ( .D(n2521), .CK(n993), .QN(lo_out[26]) );
  DFF_X1 \lo/q_reg[27]  ( .D(n2520), .CK(n993), .QN(lo_out[27]) );
  DFF_X1 \lo/q_reg[28]  ( .D(n2519), .CK(n993), .QN(lo_out[28]) );
  DFF_X1 \lo/q_reg[29]  ( .D(n2518), .CK(n993), .QN(lo_out[29]) );
  DFF_X1 \lo/q_reg[30]  ( .D(n2517), .CK(n993), .QN(lo_out[30]) );
  DFF_X1 \lo/q_reg[31]  ( .D(n2516), .CK(n993), .QN(lo_out[31]) );
  DFF_X1 \hi/q_reg[0]  ( .D(n2515), .CK(n993), .Q(n1628), .QN(hi_out[0]) );
  DFF_X1 \hi/q_reg[1]  ( .D(n2514), .CK(n993), .Q(n1651), .QN(hi_out[1]) );
  DFF_X1 \hi/q_reg[2]  ( .D(n2513), .CK(n993), .Q(n1653), .QN(hi_out[2]) );
  DFF_X1 \hi/q_reg[3]  ( .D(n2512), .CK(n993), .Q(n1648), .QN(hi_out[3]) );
  DFF_X1 \hi/q_reg[4]  ( .D(n2511), .CK(n993), .Q(n1649), .QN(hi_out[4]) );
  DFF_X1 \hi/q_reg[5]  ( .D(n2510), .CK(n993), .Q(n1623), .QN(hi_out[5]) );
  DFF_X1 \hi/q_reg[6]  ( .D(n2509), .CK(n993), .Q(n1624), .QN(hi_out[6]) );
  DFF_X1 \hi/q_reg[7]  ( .D(n2508), .CK(n993), .Q(n1625), .QN(hi_out[7]) );
  DFF_X1 \hi/q_reg[8]  ( .D(n2507), .CK(n993), .Q(n1626), .QN(hi_out[8]) );
  DFF_X1 \hi/q_reg[9]  ( .D(n2506), .CK(n993), .Q(n1627), .QN(hi_out[9]) );
  DFF_X1 \hi/q_reg[10]  ( .D(n2505), .CK(n993), .Q(n1629), .QN(hi_out[10]) );
  DFF_X1 \hi/q_reg[11]  ( .D(n2504), .CK(n993), .Q(n1630), .QN(hi_out[11]) );
  DFF_X1 \hi/q_reg[12]  ( .D(n2503), .CK(n993), .Q(n1631), .QN(hi_out[12]) );
  DFF_X1 \hi/q_reg[13]  ( .D(n2502), .CK(n993), .Q(n1632), .QN(hi_out[13]) );
  DFF_X1 \hi/q_reg[14]  ( .D(n2501), .CK(n993), .Q(n1633), .QN(hi_out[14]) );
  DFF_X1 \hi/q_reg[15]  ( .D(n2500), .CK(n993), .Q(n1634), .QN(hi_out[15]) );
  DFF_X1 \hi/q_reg[16]  ( .D(n2499), .CK(n993), .Q(n1635), .QN(hi_out[16]) );
  DFF_X1 \hi/q_reg[17]  ( .D(n2498), .CK(n993), .Q(n1650), .QN(hi_out[17]) );
  DFF_X1 \hi/q_reg[18]  ( .D(n2497), .CK(n993), .Q(n1636), .QN(hi_out[18]) );
  DFF_X1 \hi/q_reg[19]  ( .D(n2496), .CK(n993), .Q(n1637), .QN(hi_out[19]) );
  DFF_X1 \hi/q_reg[20]  ( .D(n2495), .CK(n993), .Q(n1638), .QN(hi_out[20]) );
  DFF_X1 \hi/q_reg[21]  ( .D(n2494), .CK(n993), .Q(n1639), .QN(hi_out[21]) );
  DFF_X1 \hi/q_reg[22]  ( .D(n2493), .CK(n993), .Q(n1640), .QN(hi_out[22]) );
  DFF_X1 \hi/q_reg[23]  ( .D(n2492), .CK(n993), .Q(n1641), .QN(hi_out[23]) );
  DFF_X1 \hi/q_reg[24]  ( .D(n2491), .CK(n993), .Q(n1642), .QN(hi_out[24]) );
  DFF_X1 \hi/q_reg[25]  ( .D(n2490), .CK(n993), .Q(n1652), .QN(hi_out[25]) );
  DFF_X1 \hi/q_reg[26]  ( .D(n2489), .CK(n993), .Q(n1643), .QN(hi_out[26]) );
  DFF_X1 \hi/q_reg[27]  ( .D(n2488), .CK(n993), .Q(n1644), .QN(hi_out[27]) );
  DFF_X1 \hi/q_reg[28]  ( .D(n2487), .CK(n993), .Q(n1645), .QN(hi_out[28]) );
  DFF_X1 \hi/q_reg[29]  ( .D(n2486), .CK(n993), .Q(n1646), .QN(hi_out[29]) );
  DFF_X1 \hi/q_reg[30]  ( .D(n2485), .CK(n993), .Q(n1654), .QN(hi_out[30]) );
  DFF_X1 \hi/q_reg[31]  ( .D(n2482), .CK(n993), .Q(n1647), .QN(hi_out[31]) );
  OAI22_X1 U3 ( .A1(n855), .A2(n2261), .B1(n503), .B2(n2259), .ZN(n994) );
  OAI22_X1 U4 ( .A1(n311), .A2(n2280), .B1(n55), .B2(n2255), .ZN(n995) );
  OAI22_X1 U5 ( .A1(n663), .A2(n2278), .B1(n375), .B2(n2260), .ZN(n996) );
  OAI22_X1 U6 ( .A1(n983), .A2(n2258), .B1(n407), .B2(n2270), .ZN(n997) );
  NOR4_X1 U7 ( .A1(n994), .A2(n995), .A3(n996), .A4(n997), .ZN(n998) );
  OAI22_X1 U8 ( .A1(n87), .A2(n2251), .B1(n727), .B2(n2269), .ZN(n999) );
  OAI22_X1 U9 ( .A1(n759), .A2(n2276), .B1(n23), .B2(n2264), .ZN(n1000) );
  OAI22_X1 U10 ( .A1(n247), .A2(n2263), .B1(n183), .B2(n2257), .ZN(n1001) );
  OAI22_X1 U11 ( .A1(n887), .A2(n2275), .B1(n567), .B2(n2265), .ZN(n1002) );
  NOR4_X1 U12 ( .A1(n999), .A2(n1000), .A3(n1001), .A4(n1002), .ZN(n1003) );
  OAI222_X1 U13 ( .A1(n439), .A2(n2267), .B1(n791), .B2(n2279), .C1(n471), 
        .C2(n2268), .ZN(n1004) );
  OAI22_X1 U14 ( .A1(n215), .A2(n2266), .B1(n599), .B2(n2250), .ZN(n1005) );
  OAI22_X1 U15 ( .A1(n951), .A2(n2277), .B1(n535), .B2(n2253), .ZN(n1006) );
  NOR3_X1 U16 ( .A1(n1004), .A2(n1005), .A3(n1006), .ZN(n1007) );
  OAI22_X1 U17 ( .A1(n823), .A2(n2273), .B1(n695), .B2(n2262), .ZN(n1008) );
  OAI22_X1 U18 ( .A1(n919), .A2(n2272), .B1(n343), .B2(n2256), .ZN(n1009) );
  OAI22_X1 U19 ( .A1(n119), .A2(n2274), .B1(n631), .B2(n2271), .ZN(n1010) );
  OAI22_X1 U20 ( .A1(n279), .A2(n2252), .B1(n151), .B2(n1677), .ZN(n1011) );
  NOR4_X1 U21 ( .A1(n1008), .A2(n1009), .A3(n1010), .A4(n1011), .ZN(n1012) );
  NAND4_X1 U22 ( .A1(n998), .A2(n1003), .A3(n1007), .A4(n1012), .ZN(n1013) );
  AOI22_X1 U23 ( .A1(lo_out[22]), .A2(n1679), .B1(n2282), .B2(n1013), .ZN(
        n1014) );
  OAI21_X1 U24 ( .B1(n2283), .B2(n1640), .A(n1014), .ZN(rp1[22]) );
  OAI22_X1 U25 ( .A1(n176), .A2(n3761), .B1(n624), .B2(n3755), .ZN(n1015) );
  OAI22_X1 U26 ( .A1(n560), .A2(n3782), .B1(n592), .B2(n3759), .ZN(n1016) );
  OAI22_X1 U27 ( .A1(n880), .A2(n3778), .B1(n112), .B2(n3774), .ZN(n1017) );
  OAI22_X1 U28 ( .A1(n80), .A2(n3763), .B1(n752), .B2(n3768), .ZN(n1018) );
  NOR4_X1 U29 ( .A1(n1015), .A2(n1016), .A3(n1017), .A4(n1018), .ZN(n1019) );
  OAI22_X1 U30 ( .A1(n976), .A2(n3771), .B1(n656), .B2(n3756), .ZN(n1020) );
  OAI22_X1 U31 ( .A1(n784), .A2(n3772), .B1(n432), .B2(n3760), .ZN(n1021) );
  OAI22_X1 U32 ( .A1(n496), .A2(n3757), .B1(n336), .B2(n3777), .ZN(n1022) );
  OAI22_X1 U33 ( .A1(n912), .A2(n3783), .B1(n816), .B2(n3754), .ZN(n1023) );
  NOR4_X1 U34 ( .A1(n1020), .A2(n1021), .A3(n1022), .A4(n1023), .ZN(n1024) );
  OAI222_X1 U35 ( .A1(n528), .A2(n3779), .B1(n240), .B2(n3781), .C1(n464), 
        .C2(n3766), .ZN(n1025) );
  OAI22_X1 U36 ( .A1(n304), .A2(n3764), .B1(n208), .B2(n3758), .ZN(n1026) );
  OAI22_X1 U37 ( .A1(n144), .A2(n3769), .B1(n48), .B2(n3773), .ZN(n1027) );
  NOR3_X1 U38 ( .A1(n1025), .A2(n1026), .A3(n1027), .ZN(n1028) );
  OAI22_X1 U39 ( .A1(n720), .A2(n3762), .B1(n688), .B2(n3765), .ZN(n1029) );
  OAI22_X1 U40 ( .A1(n16), .A2(n3770), .B1(n400), .B2(n3780), .ZN(n1030) );
  OAI22_X1 U41 ( .A1(n368), .A2(n3776), .B1(n272), .B2(n3775), .ZN(n1031) );
  OAI22_X1 U42 ( .A1(n848), .A2(n3767), .B1(n944), .B2(n3784), .ZN(n1032) );
  NOR4_X1 U43 ( .A1(n1029), .A2(n1030), .A3(n1031), .A4(n1032), .ZN(n1033) );
  NAND4_X1 U44 ( .A1(n1019), .A2(n1024), .A3(n1028), .A4(n1033), .ZN(n1034) );
  AOI22_X1 U45 ( .A1(lo_out[15]), .A2(n1685), .B1(n3785), .B2(n1034), .ZN(
        n1035) );
  OAI21_X1 U46 ( .B1(n1634), .B2(n3787), .A(n1035), .ZN(rp2[15]) );
  OAI22_X1 U47 ( .A1(n854), .A2(n2261), .B1(n694), .B2(n2262), .ZN(n1036) );
  OAI22_X1 U48 ( .A1(n214), .A2(n2266), .B1(n438), .B2(n2267), .ZN(n1037) );
  OAI22_X1 U49 ( .A1(n950), .A2(n2277), .B1(n758), .B2(n2276), .ZN(n1038) );
  OAI22_X1 U50 ( .A1(n598), .A2(n2250), .B1(n150), .B2(n1677), .ZN(n1039) );
  NOR4_X1 U51 ( .A1(n1036), .A2(n1037), .A3(n1038), .A4(n1039), .ZN(n1040) );
  OAI22_X1 U52 ( .A1(n918), .A2(n2272), .B1(n374), .B2(n2260), .ZN(n1041) );
  OAI22_X1 U53 ( .A1(n86), .A2(n2251), .B1(n790), .B2(n2279), .ZN(n1042) );
  OAI22_X1 U54 ( .A1(n470), .A2(n2268), .B1(n502), .B2(n2259), .ZN(n1043) );
  OAI22_X1 U55 ( .A1(n22), .A2(n2264), .B1(n310), .B2(n2280), .ZN(n1044) );
  NOR4_X1 U56 ( .A1(n1041), .A2(n1042), .A3(n1043), .A4(n1044), .ZN(n1045) );
  OAI222_X1 U57 ( .A1(n566), .A2(n2265), .B1(n726), .B2(n2269), .C1(n406), 
        .C2(n2270), .ZN(n1046) );
  OAI22_X1 U58 ( .A1(n982), .A2(n2258), .B1(n342), .B2(n2256), .ZN(n1047) );
  OAI22_X1 U59 ( .A1(n118), .A2(n2274), .B1(n278), .B2(n2252), .ZN(n1048) );
  NOR3_X1 U60 ( .A1(n1046), .A2(n1047), .A3(n1048), .ZN(n1049) );
  OAI22_X1 U61 ( .A1(n246), .A2(n2263), .B1(n630), .B2(n2271), .ZN(n1050) );
  OAI22_X1 U62 ( .A1(n182), .A2(n2257), .B1(n54), .B2(n2255), .ZN(n1051) );
  OAI22_X1 U63 ( .A1(n534), .A2(n2253), .B1(n662), .B2(n2278), .ZN(n1052) );
  OAI22_X1 U64 ( .A1(n886), .A2(n2275), .B1(n822), .B2(n2273), .ZN(n1053) );
  NOR4_X1 U65 ( .A1(n1050), .A2(n1051), .A3(n1052), .A4(n1053), .ZN(n1054) );
  NAND4_X1 U66 ( .A1(n1040), .A2(n1045), .A3(n1049), .A4(n1054), .ZN(n1055) );
  AOI22_X1 U67 ( .A1(lo_out[21]), .A2(n2281), .B1(n2282), .B2(n1055), .ZN(
        n1056) );
  OAI21_X1 U68 ( .B1(n2283), .B2(n1639), .A(n1056), .ZN(rp1[21]) );
  OAI22_X1 U69 ( .A1(n911), .A2(n3783), .B1(n335), .B2(n3777), .ZN(n1057) );
  OAI22_X1 U70 ( .A1(n463), .A2(n3766), .B1(n15), .B2(n3770), .ZN(n1058) );
  OAI22_X1 U71 ( .A1(n879), .A2(n3778), .B1(n367), .B2(n3776), .ZN(n1059) );
  OAI22_X1 U72 ( .A1(n975), .A2(n3771), .B1(n719), .B2(n3762), .ZN(n1060) );
  NOR4_X1 U73 ( .A1(n1057), .A2(n1058), .A3(n1059), .A4(n1060), .ZN(n1061) );
  OAI22_X1 U74 ( .A1(n847), .A2(n3767), .B1(n527), .B2(n3779), .ZN(n1062) );
  OAI22_X1 U75 ( .A1(n943), .A2(n3784), .B1(n751), .B2(n3768), .ZN(n1063) );
  OAI22_X1 U76 ( .A1(n175), .A2(n3761), .B1(n239), .B2(n3781), .ZN(n1064) );
  OAI22_X1 U77 ( .A1(n431), .A2(n3760), .B1(n271), .B2(n3775), .ZN(n1065) );
  NOR4_X1 U78 ( .A1(n1062), .A2(n1063), .A3(n1064), .A4(n1065), .ZN(n1066) );
  OAI222_X1 U79 ( .A1(n111), .A2(n3774), .B1(n623), .B2(n3755), .C1(n655), 
        .C2(n3756), .ZN(n1067) );
  OAI22_X1 U80 ( .A1(n591), .A2(n3759), .B1(n303), .B2(n3764), .ZN(n1068) );
  OAI22_X1 U81 ( .A1(n687), .A2(n3765), .B1(n79), .B2(n3763), .ZN(n1069) );
  NOR3_X1 U82 ( .A1(n1067), .A2(n1068), .A3(n1069), .ZN(n1070) );
  OAI22_X1 U83 ( .A1(n399), .A2(n3780), .B1(n783), .B2(n3772), .ZN(n1071) );
  OAI22_X1 U84 ( .A1(n143), .A2(n3769), .B1(n815), .B2(n3754), .ZN(n1072) );
  OAI22_X1 U85 ( .A1(n207), .A2(n3758), .B1(n559), .B2(n3782), .ZN(n1073) );
  OAI22_X1 U86 ( .A1(n47), .A2(n3773), .B1(n495), .B2(n3757), .ZN(n1074) );
  NOR4_X1 U87 ( .A1(n1071), .A2(n1072), .A3(n1073), .A4(n1074), .ZN(n1075) );
  NAND4_X1 U88 ( .A1(n1061), .A2(n1066), .A3(n1070), .A4(n1075), .ZN(n1076) );
  AOI22_X1 U89 ( .A1(lo_out[14]), .A2(n1685), .B1(n1684), .B2(n1076), .ZN(
        n1077) );
  OAI21_X1 U90 ( .B1(n1633), .B2(n3787), .A(n1077), .ZN(rp2[14]) );
  OAI22_X1 U91 ( .A1(n885), .A2(n2275), .B1(n565), .B2(n2265), .ZN(n1078) );
  OAI22_X1 U92 ( .A1(n981), .A2(n2258), .B1(n149), .B2(n2254), .ZN(n1079) );
  OAI22_X1 U93 ( .A1(n277), .A2(n2252), .B1(n661), .B2(n2278), .ZN(n1080) );
  OAI22_X1 U94 ( .A1(n693), .A2(n2262), .B1(n85), .B2(n2251), .ZN(n1081) );
  NOR4_X1 U95 ( .A1(n1078), .A2(n1079), .A3(n1080), .A4(n1081), .ZN(n1082) );
  OAI22_X1 U96 ( .A1(n213), .A2(n2266), .B1(n21), .B2(n2264), .ZN(n1083) );
  OAI22_X1 U97 ( .A1(n917), .A2(n2272), .B1(n469), .B2(n2268), .ZN(n1084) );
  OAI22_X1 U98 ( .A1(n949), .A2(n2277), .B1(n373), .B2(n2260), .ZN(n1085) );
  OAI22_X1 U99 ( .A1(n245), .A2(n2263), .B1(n181), .B2(n2257), .ZN(n1086) );
  NOR4_X1 U100 ( .A1(n1083), .A2(n1084), .A3(n1085), .A4(n1086), .ZN(n1087) );
  OAI222_X1 U101 ( .A1(n629), .A2(n2271), .B1(n789), .B2(n2279), .C1(n309), 
        .C2(n2280), .ZN(n1088) );
  OAI22_X1 U102 ( .A1(n53), .A2(n2255), .B1(n725), .B2(n2269), .ZN(n1089) );
  OAI22_X1 U103 ( .A1(n533), .A2(n2253), .B1(n117), .B2(n2274), .ZN(n1090) );
  NOR3_X1 U104 ( .A1(n1088), .A2(n1089), .A3(n1090), .ZN(n1091) );
  OAI22_X1 U105 ( .A1(n405), .A2(n2270), .B1(n757), .B2(n2276), .ZN(n1092) );
  OAI22_X1 U106 ( .A1(n597), .A2(n2250), .B1(n501), .B2(n2259), .ZN(n1093) );
  OAI22_X1 U107 ( .A1(n853), .A2(n2261), .B1(n437), .B2(n2267), .ZN(n1094) );
  OAI22_X1 U108 ( .A1(n341), .A2(n2256), .B1(n821), .B2(n2273), .ZN(n1095) );
  NOR4_X1 U109 ( .A1(n1092), .A2(n1093), .A3(n1094), .A4(n1095), .ZN(n1096) );
  NAND4_X1 U110 ( .A1(n1082), .A2(n1087), .A3(n1091), .A4(n1096), .ZN(n1097)
         );
  AOI22_X1 U111 ( .A1(lo_out[20]), .A2(n1679), .B1(n2282), .B2(n1097), .ZN(
        n1098) );
  OAI21_X1 U112 ( .B1(n2283), .B2(n1638), .A(n1098), .ZN(rp1[20]) );
  OAI22_X1 U113 ( .A1(n878), .A2(n3778), .B1(n462), .B2(n3766), .ZN(n1099) );
  OAI22_X1 U114 ( .A1(n238), .A2(n3781), .B1(n558), .B2(n3782), .ZN(n1100) );
  OAI22_X1 U115 ( .A1(n270), .A2(n3775), .B1(n398), .B2(n1683), .ZN(n1101) );
  OAI22_X1 U116 ( .A1(n206), .A2(n3758), .B1(n654), .B2(n3756), .ZN(n1102) );
  NOR4_X1 U117 ( .A1(n1099), .A2(n1100), .A3(n1101), .A4(n1102), .ZN(n1103) );
  OAI22_X1 U118 ( .A1(n782), .A2(n3772), .B1(n526), .B2(n3779), .ZN(n1104) );
  OAI22_X1 U119 ( .A1(n750), .A2(n3768), .B1(n430), .B2(n3760), .ZN(n1105) );
  OAI22_X1 U120 ( .A1(n814), .A2(n3754), .B1(n590), .B2(n3759), .ZN(n1106) );
  OAI22_X1 U121 ( .A1(n846), .A2(n3767), .B1(n974), .B2(n3771), .ZN(n1107) );
  NOR4_X1 U122 ( .A1(n1104), .A2(n1105), .A3(n1106), .A4(n1107), .ZN(n1108) );
  OAI222_X1 U123 ( .A1(n686), .A2(n3765), .B1(n366), .B2(n3776), .C1(n334), 
        .C2(n3777), .ZN(n1109) );
  OAI22_X1 U124 ( .A1(n302), .A2(n3764), .B1(n174), .B2(n3761), .ZN(n1110) );
  OAI22_X1 U125 ( .A1(n110), .A2(n3774), .B1(n142), .B2(n3769), .ZN(n1111) );
  NOR3_X1 U126 ( .A1(n1109), .A2(n1110), .A3(n1111), .ZN(n1112) );
  OAI22_X1 U127 ( .A1(n718), .A2(n3762), .B1(n14), .B2(n3770), .ZN(n1113) );
  OAI22_X1 U128 ( .A1(n622), .A2(n1681), .B1(n494), .B2(n3757), .ZN(n1114) );
  OAI22_X1 U129 ( .A1(n910), .A2(n3783), .B1(n78), .B2(n3763), .ZN(n1115) );
  OAI22_X1 U130 ( .A1(n942), .A2(n3784), .B1(n46), .B2(n3773), .ZN(n1116) );
  NOR4_X1 U131 ( .A1(n1113), .A2(n1114), .A3(n1115), .A4(n1116), .ZN(n1117) );
  NAND4_X1 U132 ( .A1(n1103), .A2(n1108), .A3(n1112), .A4(n1117), .ZN(n1118)
         );
  AOI22_X1 U133 ( .A1(lo_out[13]), .A2(n1685), .B1(n3785), .B2(n1118), .ZN(
        n1119) );
  OAI21_X1 U134 ( .B1(n1632), .B2(n3787), .A(n1119), .ZN(rp2[13]) );
  OAI22_X1 U135 ( .A1(n300), .A2(n2280), .B1(n780), .B2(n2279), .ZN(n1120) );
  OAI22_X1 U136 ( .A1(n396), .A2(n2270), .B1(n108), .B2(n2274), .ZN(n1121) );
  OAI22_X1 U137 ( .A1(n204), .A2(n2266), .B1(n844), .B2(n2261), .ZN(n1122) );
  OAI22_X1 U138 ( .A1(n12), .A2(n2264), .B1(n812), .B2(n2273), .ZN(n1123) );
  NOR4_X1 U139 ( .A1(n1120), .A2(n1121), .A3(n1122), .A4(n1123), .ZN(n1124) );
  OAI22_X1 U140 ( .A1(n908), .A2(n2272), .B1(n716), .B2(n2269), .ZN(n1125) );
  OAI22_X1 U141 ( .A1(n492), .A2(n2259), .B1(n972), .B2(n2258), .ZN(n1126) );
  OAI22_X1 U142 ( .A1(n876), .A2(n2275), .B1(n524), .B2(n2253), .ZN(n1127) );
  OAI22_X1 U143 ( .A1(n236), .A2(n2263), .B1(n556), .B2(n2265), .ZN(n1128) );
  NOR4_X1 U144 ( .A1(n1125), .A2(n1126), .A3(n1127), .A4(n1128), .ZN(n1129) );
  OAI222_X1 U145 ( .A1(n652), .A2(n2278), .B1(n76), .B2(n2251), .C1(n172), 
        .C2(n2257), .ZN(n1130) );
  OAI22_X1 U146 ( .A1(n588), .A2(n2250), .B1(n44), .B2(n2255), .ZN(n1131) );
  OAI22_X1 U147 ( .A1(n940), .A2(n2277), .B1(n620), .B2(n1678), .ZN(n1132) );
  NOR3_X1 U148 ( .A1(n1130), .A2(n1131), .A3(n1132), .ZN(n1133) );
  OAI22_X1 U149 ( .A1(n364), .A2(n2260), .B1(n428), .B2(n2267), .ZN(n1134) );
  OAI22_X1 U150 ( .A1(n460), .A2(n2268), .B1(n140), .B2(n2254), .ZN(n1135) );
  OAI22_X1 U151 ( .A1(n332), .A2(n2256), .B1(n748), .B2(n2276), .ZN(n1136) );
  OAI22_X1 U152 ( .A1(n684), .A2(n2262), .B1(n268), .B2(n2252), .ZN(n1137) );
  NOR4_X1 U153 ( .A1(n1134), .A2(n1135), .A3(n1136), .A4(n1137), .ZN(n1138) );
  NAND4_X1 U154 ( .A1(n1124), .A2(n1129), .A3(n1133), .A4(n1138), .ZN(n1139)
         );
  AOI22_X1 U155 ( .A1(lo_out[11]), .A2(n1679), .B1(n2282), .B2(n1139), .ZN(
        n1140) );
  OAI21_X1 U156 ( .B1(n2283), .B2(n1630), .A(n1140), .ZN(rp1[11]) );
  OAI22_X1 U157 ( .A1(n237), .A2(n3781), .B1(n813), .B2(n3754), .ZN(n1141) );
  OAI22_X1 U158 ( .A1(n941), .A2(n3784), .B1(n301), .B2(n3764), .ZN(n1142) );
  OAI22_X1 U159 ( .A1(n173), .A2(n3761), .B1(n845), .B2(n3767), .ZN(n1143) );
  OAI22_X1 U160 ( .A1(n717), .A2(n3762), .B1(n333), .B2(n3777), .ZN(n1144) );
  NOR4_X1 U161 ( .A1(n1141), .A2(n1142), .A3(n1143), .A4(n1144), .ZN(n1145) );
  OAI22_X1 U162 ( .A1(n653), .A2(n3756), .B1(n557), .B2(n3782), .ZN(n1146) );
  OAI22_X1 U163 ( .A1(n13), .A2(n3770), .B1(n77), .B2(n3763), .ZN(n1147) );
  OAI22_X1 U164 ( .A1(n429), .A2(n3760), .B1(n461), .B2(n3766), .ZN(n1148) );
  OAI22_X1 U165 ( .A1(n621), .A2(n3755), .B1(n365), .B2(n3776), .ZN(n1149) );
  NOR4_X1 U166 ( .A1(n1146), .A2(n1147), .A3(n1148), .A4(n1149), .ZN(n1150) );
  OAI222_X1 U167 ( .A1(n205), .A2(n3758), .B1(n109), .B2(n3774), .C1(n493), 
        .C2(n3757), .ZN(n1151) );
  OAI22_X1 U168 ( .A1(n781), .A2(n3772), .B1(n141), .B2(n3769), .ZN(n1152) );
  OAI22_X1 U169 ( .A1(n749), .A2(n3768), .B1(n589), .B2(n3759), .ZN(n1153) );
  NOR3_X1 U170 ( .A1(n1151), .A2(n1152), .A3(n1153), .ZN(n1154) );
  OAI22_X1 U171 ( .A1(n525), .A2(n3779), .B1(n973), .B2(n3771), .ZN(n1155) );
  OAI22_X1 U172 ( .A1(n45), .A2(n3773), .B1(n685), .B2(n3765), .ZN(n1156) );
  OAI22_X1 U173 ( .A1(n877), .A2(n3778), .B1(n269), .B2(n3775), .ZN(n1157) );
  OAI22_X1 U174 ( .A1(n909), .A2(n3783), .B1(n397), .B2(n3780), .ZN(n1158) );
  NOR4_X1 U175 ( .A1(n1155), .A2(n1156), .A3(n1157), .A4(n1158), .ZN(n1159) );
  NAND4_X1 U176 ( .A1(n1145), .A2(n1150), .A3(n1154), .A4(n1159), .ZN(n1160)
         );
  AOI22_X1 U177 ( .A1(lo_out[12]), .A2(n1685), .B1(n3785), .B2(n1160), .ZN(
        n1161) );
  OAI21_X1 U178 ( .B1(n1631), .B2(n3787), .A(n1161), .ZN(rp2[12]) );
  OAI22_X1 U179 ( .A1(n148), .A2(n2254), .B1(n500), .B2(n2259), .ZN(n1162) );
  OAI22_X1 U180 ( .A1(n116), .A2(n2274), .B1(n756), .B2(n2276), .ZN(n1163) );
  OAI22_X1 U181 ( .A1(n948), .A2(n2277), .B1(n820), .B2(n2273), .ZN(n1164) );
  OAI22_X1 U182 ( .A1(n980), .A2(n2258), .B1(n308), .B2(n2280), .ZN(n1165) );
  NOR4_X1 U183 ( .A1(n1162), .A2(n1163), .A3(n1164), .A4(n1165), .ZN(n1166) );
  OAI22_X1 U184 ( .A1(n532), .A2(n2253), .B1(n692), .B2(n2262), .ZN(n1167) );
  OAI22_X1 U185 ( .A1(n916), .A2(n2272), .B1(n788), .B2(n2279), .ZN(n1168) );
  OAI22_X1 U186 ( .A1(n852), .A2(n2261), .B1(n628), .B2(n2271), .ZN(n1169) );
  OAI22_X1 U187 ( .A1(n276), .A2(n2252), .B1(n884), .B2(n2275), .ZN(n1170) );
  NOR4_X1 U188 ( .A1(n1167), .A2(n1168), .A3(n1169), .A4(n1170), .ZN(n1171) );
  OAI222_X1 U189 ( .A1(n84), .A2(n2251), .B1(n724), .B2(n2269), .C1(n180), 
        .C2(n2257), .ZN(n1172) );
  OAI22_X1 U190 ( .A1(n660), .A2(n2278), .B1(n404), .B2(n2270), .ZN(n1173) );
  OAI22_X1 U191 ( .A1(n564), .A2(n2265), .B1(n468), .B2(n2268), .ZN(n1174) );
  NOR3_X1 U192 ( .A1(n1172), .A2(n1173), .A3(n1174), .ZN(n1175) );
  OAI22_X1 U193 ( .A1(n212), .A2(n2266), .B1(n340), .B2(n2256), .ZN(n1176) );
  OAI22_X1 U194 ( .A1(n244), .A2(n2263), .B1(n52), .B2(n2255), .ZN(n1177) );
  OAI22_X1 U195 ( .A1(n596), .A2(n2250), .B1(n372), .B2(n2260), .ZN(n1178) );
  OAI22_X1 U196 ( .A1(n20), .A2(n2264), .B1(n436), .B2(n2267), .ZN(n1179) );
  NOR4_X1 U197 ( .A1(n1176), .A2(n1177), .A3(n1178), .A4(n1179), .ZN(n1180) );
  NAND4_X1 U198 ( .A1(n1166), .A2(n1171), .A3(n1175), .A4(n1180), .ZN(n1181)
         );
  AOI22_X1 U199 ( .A1(lo_out[19]), .A2(n2281), .B1(n1680), .B2(n1181), .ZN(
        n1182) );
  OAI21_X1 U200 ( .B1(n2283), .B2(n1637), .A(n1182), .ZN(rp1[19]) );
  OAI22_X1 U201 ( .A1(n12), .A2(n3770), .B1(n492), .B2(n3757), .ZN(n1183) );
  OAI22_X1 U202 ( .A1(n940), .A2(n3784), .B1(n652), .B2(n3756), .ZN(n1184) );
  OAI22_X1 U203 ( .A1(n204), .A2(n3758), .B1(n780), .B2(n3772), .ZN(n1185) );
  OAI22_X1 U204 ( .A1(n972), .A2(n3771), .B1(n908), .B2(n3783), .ZN(n1186) );
  NOR4_X1 U205 ( .A1(n1183), .A2(n1184), .A3(n1185), .A4(n1186), .ZN(n1187) );
  OAI22_X1 U206 ( .A1(n332), .A2(n3777), .B1(n140), .B2(n3769), .ZN(n1188) );
  OAI22_X1 U207 ( .A1(n716), .A2(n3762), .B1(n556), .B2(n3782), .ZN(n1189) );
  OAI22_X1 U208 ( .A1(n108), .A2(n3774), .B1(n396), .B2(n3780), .ZN(n1190) );
  OAI22_X1 U209 ( .A1(n300), .A2(n3764), .B1(n588), .B2(n3759), .ZN(n1191) );
  NOR4_X1 U210 ( .A1(n1188), .A2(n1189), .A3(n1190), .A4(n1191), .ZN(n1192) );
  OAI222_X1 U211 ( .A1(n876), .A2(n3778), .B1(n812), .B2(n3754), .C1(n748), 
        .C2(n3768), .ZN(n1193) );
  OAI22_X1 U212 ( .A1(n76), .A2(n3763), .B1(n428), .B2(n3760), .ZN(n1194) );
  OAI22_X1 U213 ( .A1(n172), .A2(n3761), .B1(n44), .B2(n3773), .ZN(n1195) );
  NOR3_X1 U214 ( .A1(n1193), .A2(n1194), .A3(n1195), .ZN(n1196) );
  OAI22_X1 U215 ( .A1(n460), .A2(n3766), .B1(n364), .B2(n3776), .ZN(n1197) );
  OAI22_X1 U216 ( .A1(n844), .A2(n3767), .B1(n524), .B2(n3779), .ZN(n1198) );
  OAI22_X1 U217 ( .A1(n268), .A2(n3775), .B1(n620), .B2(n1681), .ZN(n1199) );
  OAI22_X1 U218 ( .A1(n684), .A2(n3765), .B1(n236), .B2(n3781), .ZN(n1200) );
  NOR4_X1 U219 ( .A1(n1197), .A2(n1198), .A3(n1199), .A4(n1200), .ZN(n1201) );
  NAND4_X1 U220 ( .A1(n1187), .A2(n1192), .A3(n1196), .A4(n1201), .ZN(n1202)
         );
  AOI22_X1 U221 ( .A1(lo_out[11]), .A2(n1685), .B1(n1684), .B2(n1202), .ZN(
        n1203) );
  OAI21_X1 U222 ( .B1(n1630), .B2(n3787), .A(n1203), .ZN(rp2[11]) );
  OAI22_X1 U223 ( .A1(n554), .A2(n2265), .B1(n202), .B2(n2266), .ZN(n1204) );
  OAI22_X1 U224 ( .A1(n426), .A2(n2267), .B1(n458), .B2(n2268), .ZN(n1205) );
  OAI22_X1 U225 ( .A1(n714), .A2(n2269), .B1(n394), .B2(n2270), .ZN(n1206) );
  OAI22_X1 U226 ( .A1(n618), .A2(n1678), .B1(n906), .B2(n2272), .ZN(n1207) );
  NOR4_X1 U227 ( .A1(n1204), .A2(n1205), .A3(n1206), .A4(n1207), .ZN(n1208) );
  OAI22_X1 U228 ( .A1(n810), .A2(n2273), .B1(n106), .B2(n2274), .ZN(n1209) );
  OAI22_X1 U229 ( .A1(n874), .A2(n2275), .B1(n746), .B2(n2276), .ZN(n1210) );
  OAI22_X1 U230 ( .A1(n938), .A2(n2277), .B1(n650), .B2(n2278), .ZN(n1211) );
  OAI22_X1 U231 ( .A1(n778), .A2(n2279), .B1(n298), .B2(n2280), .ZN(n1212) );
  NOR4_X1 U232 ( .A1(n1209), .A2(n1210), .A3(n1211), .A4(n1212), .ZN(n1213) );
  OAI222_X1 U233 ( .A1(n74), .A2(n2251), .B1(n266), .B2(n2252), .C1(n586), 
        .C2(n2250), .ZN(n1214) );
  OAI22_X1 U234 ( .A1(n522), .A2(n2253), .B1(n138), .B2(n1677), .ZN(n1215) );
  OAI22_X1 U235 ( .A1(n42), .A2(n2255), .B1(n330), .B2(n2256), .ZN(n1216) );
  NOR3_X1 U236 ( .A1(n1214), .A2(n1215), .A3(n1216), .ZN(n1217) );
  OAI22_X1 U237 ( .A1(n170), .A2(n2257), .B1(n970), .B2(n2258), .ZN(n1218) );
  OAI22_X1 U238 ( .A1(n490), .A2(n2259), .B1(n362), .B2(n2260), .ZN(n1219) );
  OAI22_X1 U239 ( .A1(n842), .A2(n2261), .B1(n682), .B2(n2262), .ZN(n1220) );
  OAI22_X1 U240 ( .A1(n234), .A2(n2263), .B1(n10), .B2(n2264), .ZN(n1221) );
  NOR4_X1 U241 ( .A1(n1218), .A2(n1219), .A3(n1220), .A4(n1221), .ZN(n1222) );
  NAND4_X1 U242 ( .A1(n1208), .A2(n1213), .A3(n1217), .A4(n1222), .ZN(n1223)
         );
  AOI22_X1 U243 ( .A1(lo_out[9]), .A2(n1679), .B1(n1680), .B2(n1223), .ZN(
        n1224) );
  OAI21_X1 U244 ( .B1(n2283), .B2(n1627), .A(n1224), .ZN(rp1[9]) );
  OAI22_X1 U245 ( .A1(n555), .A2(n3782), .B1(n971), .B2(n3771), .ZN(n1225) );
  OAI22_X1 U246 ( .A1(n331), .A2(n3777), .B1(n395), .B2(n1683), .ZN(n1226) );
  OAI22_X1 U247 ( .A1(n43), .A2(n3773), .B1(n715), .B2(n3762), .ZN(n1227) );
  OAI22_X1 U248 ( .A1(n427), .A2(n3760), .B1(n299), .B2(n3764), .ZN(n1228) );
  NOR4_X1 U249 ( .A1(n1225), .A2(n1226), .A3(n1227), .A4(n1228), .ZN(n1229) );
  OAI22_X1 U250 ( .A1(n587), .A2(n3759), .B1(n843), .B2(n3767), .ZN(n1230) );
  OAI22_X1 U251 ( .A1(n875), .A2(n3778), .B1(n363), .B2(n3776), .ZN(n1231) );
  OAI22_X1 U252 ( .A1(n651), .A2(n3756), .B1(n907), .B2(n3783), .ZN(n1232) );
  OAI22_X1 U253 ( .A1(n491), .A2(n3757), .B1(n235), .B2(n3781), .ZN(n1233) );
  NOR4_X1 U254 ( .A1(n1230), .A2(n1231), .A3(n1232), .A4(n1233), .ZN(n1234) );
  OAI222_X1 U255 ( .A1(n619), .A2(n3755), .B1(n779), .B2(n3772), .C1(n107), 
        .C2(n3774), .ZN(n1235) );
  OAI22_X1 U256 ( .A1(n267), .A2(n3775), .B1(n811), .B2(n3754), .ZN(n1236) );
  OAI22_X1 U257 ( .A1(n11), .A2(n3770), .B1(n459), .B2(n3766), .ZN(n1237) );
  NOR3_X1 U258 ( .A1(n1235), .A2(n1236), .A3(n1237), .ZN(n1238) );
  OAI22_X1 U259 ( .A1(n523), .A2(n3779), .B1(n683), .B2(n3765), .ZN(n1239) );
  OAI22_X1 U260 ( .A1(n939), .A2(n3784), .B1(n75), .B2(n3763), .ZN(n1240) );
  OAI22_X1 U261 ( .A1(n203), .A2(n3758), .B1(n171), .B2(n3761), .ZN(n1241) );
  OAI22_X1 U262 ( .A1(n747), .A2(n3768), .B1(n139), .B2(n3769), .ZN(n1242) );
  NOR4_X1 U263 ( .A1(n1239), .A2(n1240), .A3(n1241), .A4(n1242), .ZN(n1243) );
  NAND4_X1 U264 ( .A1(n1229), .A2(n1234), .A3(n1238), .A4(n1243), .ZN(n1244)
         );
  AOI22_X1 U265 ( .A1(lo_out[10]), .A2(n1685), .B1(n1684), .B2(n1244), .ZN(
        n1245) );
  OAI21_X1 U266 ( .B1(n1629), .B2(n3787), .A(n1245), .ZN(rp2[10]) );
  OAI22_X1 U267 ( .A1(n173), .A2(n2257), .B1(n525), .B2(n2253), .ZN(n1246) );
  OAI22_X1 U268 ( .A1(n653), .A2(n2278), .B1(n781), .B2(n2279), .ZN(n1247) );
  OAI22_X1 U269 ( .A1(n909), .A2(n2272), .B1(n589), .B2(n2250), .ZN(n1248) );
  OAI22_X1 U270 ( .A1(n493), .A2(n2259), .B1(n429), .B2(n2267), .ZN(n1249) );
  NOR4_X1 U271 ( .A1(n1246), .A2(n1247), .A3(n1248), .A4(n1249), .ZN(n1250) );
  OAI22_X1 U272 ( .A1(n237), .A2(n2263), .B1(n877), .B2(n2275), .ZN(n1251) );
  OAI22_X1 U273 ( .A1(n461), .A2(n2268), .B1(n77), .B2(n2251), .ZN(n1252) );
  OAI22_X1 U274 ( .A1(n397), .A2(n2270), .B1(n109), .B2(n2274), .ZN(n1253) );
  OAI22_X1 U275 ( .A1(n813), .A2(n2273), .B1(n141), .B2(n2254), .ZN(n1254) );
  NOR4_X1 U276 ( .A1(n1251), .A2(n1252), .A3(n1253), .A4(n1254), .ZN(n1255) );
  OAI222_X1 U277 ( .A1(n717), .A2(n2269), .B1(n845), .B2(n2261), .C1(n333), 
        .C2(n2256), .ZN(n1256) );
  OAI22_X1 U278 ( .A1(n45), .A2(n2255), .B1(n13), .B2(n2264), .ZN(n1257) );
  OAI22_X1 U279 ( .A1(n205), .A2(n2266), .B1(n301), .B2(n2280), .ZN(n1258) );
  NOR3_X1 U280 ( .A1(n1256), .A2(n1257), .A3(n1258), .ZN(n1259) );
  OAI22_X1 U281 ( .A1(n749), .A2(n2276), .B1(n269), .B2(n2252), .ZN(n1260) );
  OAI22_X1 U282 ( .A1(n941), .A2(n2277), .B1(n365), .B2(n2260), .ZN(n1261) );
  OAI22_X1 U283 ( .A1(n973), .A2(n2258), .B1(n685), .B2(n2262), .ZN(n1262) );
  OAI22_X1 U284 ( .A1(n621), .A2(n1678), .B1(n557), .B2(n2265), .ZN(n1263) );
  NOR4_X1 U285 ( .A1(n1260), .A2(n1261), .A3(n1262), .A4(n1263), .ZN(n1264) );
  NAND4_X1 U286 ( .A1(n1250), .A2(n1255), .A3(n1259), .A4(n1264), .ZN(n1265)
         );
  AOI22_X1 U287 ( .A1(lo_out[12]), .A2(n1679), .B1(n2282), .B2(n1265), .ZN(
        n1266) );
  OAI21_X1 U288 ( .B1(n2283), .B2(n1631), .A(n1266), .ZN(rp1[12]) );
  OAI22_X1 U289 ( .A1(n138), .A2(n1682), .B1(n10), .B2(n3770), .ZN(n1267) );
  OAI22_X1 U290 ( .A1(n778), .A2(n3772), .B1(n970), .B2(n3771), .ZN(n1268) );
  OAI22_X1 U291 ( .A1(n106), .A2(n3774), .B1(n42), .B2(n3773), .ZN(n1269) );
  OAI22_X1 U292 ( .A1(n362), .A2(n3776), .B1(n266), .B2(n3775), .ZN(n1270) );
  NOR4_X1 U293 ( .A1(n1267), .A2(n1268), .A3(n1269), .A4(n1270), .ZN(n1271) );
  OAI22_X1 U294 ( .A1(n874), .A2(n3778), .B1(n330), .B2(n3777), .ZN(n1272) );
  OAI22_X1 U295 ( .A1(n522), .A2(n3779), .B1(n394), .B2(n3780), .ZN(n1273) );
  OAI22_X1 U296 ( .A1(n234), .A2(n3781), .B1(n554), .B2(n3782), .ZN(n1274) );
  OAI22_X1 U297 ( .A1(n938), .A2(n3784), .B1(n906), .B2(n3783), .ZN(n1275) );
  NOR4_X1 U298 ( .A1(n1272), .A2(n1273), .A3(n1274), .A4(n1275), .ZN(n1276) );
  OAI222_X1 U299 ( .A1(n810), .A2(n3754), .B1(n650), .B2(n3756), .C1(n618), 
        .C2(n1681), .ZN(n1277) );
  OAI22_X1 U300 ( .A1(n490), .A2(n3757), .B1(n202), .B2(n3758), .ZN(n1278) );
  OAI22_X1 U301 ( .A1(n586), .A2(n3759), .B1(n426), .B2(n3760), .ZN(n1279) );
  NOR3_X1 U302 ( .A1(n1277), .A2(n1278), .A3(n1279), .ZN(n1280) );
  OAI22_X1 U303 ( .A1(n714), .A2(n3762), .B1(n170), .B2(n3761), .ZN(n1281) );
  OAI22_X1 U304 ( .A1(n74), .A2(n3763), .B1(n298), .B2(n3764), .ZN(n1282) );
  OAI22_X1 U305 ( .A1(n458), .A2(n3766), .B1(n682), .B2(n3765), .ZN(n1283) );
  OAI22_X1 U306 ( .A1(n842), .A2(n3767), .B1(n746), .B2(n3768), .ZN(n1284) );
  NOR4_X1 U307 ( .A1(n1281), .A2(n1282), .A3(n1283), .A4(n1284), .ZN(n1285) );
  NAND4_X1 U308 ( .A1(n1271), .A2(n1276), .A3(n1280), .A4(n1285), .ZN(n1286)
         );
  AOI22_X1 U309 ( .A1(lo_out[9]), .A2(n3786), .B1(n1684), .B2(n1286), .ZN(
        n1287) );
  OAI21_X1 U310 ( .B1(n1627), .B2(n3787), .A(n1287), .ZN(rp2[9]) );
  OAI22_X1 U311 ( .A1(n489), .A2(n2259), .B1(n905), .B2(n2272), .ZN(n1288) );
  OAI22_X1 U312 ( .A1(n553), .A2(n2265), .B1(n937), .B2(n2277), .ZN(n1289) );
  OAI22_X1 U313 ( .A1(n841), .A2(n2261), .B1(n457), .B2(n2268), .ZN(n1290) );
  OAI22_X1 U314 ( .A1(n201), .A2(n2266), .B1(n73), .B2(n2251), .ZN(n1291) );
  NOR4_X1 U315 ( .A1(n1288), .A2(n1289), .A3(n1290), .A4(n1291), .ZN(n1292) );
  OAI22_X1 U316 ( .A1(n777), .A2(n2279), .B1(n297), .B2(n2280), .ZN(n1293) );
  OAI22_X1 U317 ( .A1(n521), .A2(n2253), .B1(n105), .B2(n2274), .ZN(n1294) );
  OAI22_X1 U318 ( .A1(n649), .A2(n2278), .B1(n9), .B2(n2264), .ZN(n1295) );
  OAI22_X1 U319 ( .A1(n265), .A2(n2252), .B1(n809), .B2(n2273), .ZN(n1296) );
  NOR4_X1 U320 ( .A1(n1293), .A2(n1294), .A3(n1295), .A4(n1296), .ZN(n1297) );
  OAI222_X1 U321 ( .A1(n713), .A2(n2269), .B1(n169), .B2(n2257), .C1(n969), 
        .C2(n2258), .ZN(n1298) );
  OAI22_X1 U322 ( .A1(n361), .A2(n2260), .B1(n585), .B2(n2250), .ZN(n1299) );
  OAI22_X1 U323 ( .A1(n425), .A2(n2267), .B1(n745), .B2(n2276), .ZN(n1300) );
  NOR3_X1 U324 ( .A1(n1298), .A2(n1299), .A3(n1300), .ZN(n1301) );
  OAI22_X1 U325 ( .A1(n393), .A2(n2270), .B1(n873), .B2(n2275), .ZN(n1302) );
  OAI22_X1 U326 ( .A1(n137), .A2(n2254), .B1(n681), .B2(n2262), .ZN(n1303) );
  OAI22_X1 U327 ( .A1(n233), .A2(n2263), .B1(n329), .B2(n2256), .ZN(n1304) );
  OAI22_X1 U328 ( .A1(n41), .A2(n2255), .B1(n617), .B2(n1678), .ZN(n1305) );
  NOR4_X1 U329 ( .A1(n1302), .A2(n1303), .A3(n1304), .A4(n1305), .ZN(n1306) );
  NAND4_X1 U330 ( .A1(n1292), .A2(n1297), .A3(n1301), .A4(n1306), .ZN(n1307)
         );
  AOI22_X1 U331 ( .A1(lo_out[8]), .A2(n1679), .B1(n1680), .B2(n1307), .ZN(
        n1308) );
  OAI21_X1 U332 ( .B1(n2283), .B2(n1626), .A(n1308), .ZN(rp1[8]) );
  OAI22_X1 U333 ( .A1(n264), .A2(n3775), .B1(n520), .B2(n3779), .ZN(n1309) );
  OAI22_X1 U334 ( .A1(n712), .A2(n3762), .B1(n136), .B2(n3769), .ZN(n1310) );
  OAI22_X1 U335 ( .A1(n200), .A2(n3758), .B1(n808), .B2(n3754), .ZN(n1311) );
  OAI22_X1 U336 ( .A1(n104), .A2(n3774), .B1(n40), .B2(n3773), .ZN(n1312) );
  NOR4_X1 U337 ( .A1(n1309), .A2(n1310), .A3(n1311), .A4(n1312), .ZN(n1313) );
  OAI22_X1 U338 ( .A1(n424), .A2(n3760), .B1(n584), .B2(n3759), .ZN(n1314) );
  OAI22_X1 U339 ( .A1(n968), .A2(n3771), .B1(n936), .B2(n3784), .ZN(n1315) );
  OAI22_X1 U340 ( .A1(n872), .A2(n3778), .B1(n296), .B2(n3764), .ZN(n1316) );
  OAI22_X1 U341 ( .A1(n616), .A2(n3755), .B1(n168), .B2(n3761), .ZN(n1317) );
  NOR4_X1 U342 ( .A1(n1314), .A2(n1315), .A3(n1316), .A4(n1317), .ZN(n1318) );
  OAI222_X1 U343 ( .A1(n328), .A2(n3777), .B1(n648), .B2(n3756), .C1(n232), 
        .C2(n3781), .ZN(n1319) );
  OAI22_X1 U344 ( .A1(n488), .A2(n3757), .B1(n776), .B2(n3772), .ZN(n1320) );
  OAI22_X1 U345 ( .A1(n744), .A2(n3768), .B1(n552), .B2(n3782), .ZN(n1321) );
  NOR3_X1 U346 ( .A1(n1319), .A2(n1320), .A3(n1321), .ZN(n1322) );
  OAI22_X1 U347 ( .A1(n392), .A2(n3780), .B1(n904), .B2(n3783), .ZN(n1323) );
  OAI22_X1 U348 ( .A1(n456), .A2(n3766), .B1(n840), .B2(n3767), .ZN(n1324) );
  OAI22_X1 U349 ( .A1(n360), .A2(n3776), .B1(n8), .B2(n3770), .ZN(n1325) );
  OAI22_X1 U350 ( .A1(n680), .A2(n3765), .B1(n72), .B2(n3763), .ZN(n1326) );
  NOR4_X1 U351 ( .A1(n1323), .A2(n1324), .A3(n1325), .A4(n1326), .ZN(n1327) );
  NAND4_X1 U352 ( .A1(n1313), .A2(n1318), .A3(n1322), .A4(n1327), .ZN(n1328)
         );
  AOI22_X1 U353 ( .A1(lo_out[7]), .A2(n3786), .B1(n1684), .B2(n1328), .ZN(
        n1329) );
  OAI21_X1 U354 ( .B1(n1625), .B2(n3787), .A(n1329), .ZN(rp2[7]) );
  OAI22_X1 U355 ( .A1(n651), .A2(n2278), .B1(n811), .B2(n2273), .ZN(n1330) );
  OAI22_X1 U356 ( .A1(n587), .A2(n2250), .B1(n683), .B2(n2262), .ZN(n1331) );
  OAI22_X1 U357 ( .A1(n523), .A2(n2253), .B1(n43), .B2(n2255), .ZN(n1332) );
  OAI22_X1 U358 ( .A1(n331), .A2(n2256), .B1(n75), .B2(n2251), .ZN(n1333) );
  NOR4_X1 U359 ( .A1(n1330), .A2(n1331), .A3(n1332), .A4(n1333), .ZN(n1334) );
  OAI22_X1 U360 ( .A1(n11), .A2(n2264), .B1(n907), .B2(n2272), .ZN(n1335) );
  OAI22_X1 U361 ( .A1(n203), .A2(n2266), .B1(n427), .B2(n2267), .ZN(n1336) );
  OAI22_X1 U362 ( .A1(n971), .A2(n2258), .B1(n459), .B2(n2268), .ZN(n1337) );
  OAI22_X1 U363 ( .A1(n139), .A2(n2254), .B1(n363), .B2(n2260), .ZN(n1338) );
  NOR4_X1 U364 ( .A1(n1335), .A2(n1336), .A3(n1337), .A4(n1338), .ZN(n1339) );
  OAI222_X1 U365 ( .A1(n107), .A2(n2274), .B1(n875), .B2(n2275), .C1(n171), 
        .C2(n2257), .ZN(n1340) );
  OAI22_X1 U366 ( .A1(n299), .A2(n2280), .B1(n939), .B2(n2277), .ZN(n1341) );
  OAI22_X1 U367 ( .A1(n267), .A2(n2252), .B1(n235), .B2(n2263), .ZN(n1342) );
  NOR3_X1 U368 ( .A1(n1340), .A2(n1341), .A3(n1342), .ZN(n1343) );
  OAI22_X1 U369 ( .A1(n747), .A2(n2276), .B1(n555), .B2(n2265), .ZN(n1344) );
  OAI22_X1 U370 ( .A1(n619), .A2(n2271), .B1(n843), .B2(n2261), .ZN(n1345) );
  OAI22_X1 U371 ( .A1(n715), .A2(n2269), .B1(n491), .B2(n2259), .ZN(n1346) );
  OAI22_X1 U372 ( .A1(n395), .A2(n2270), .B1(n779), .B2(n2279), .ZN(n1347) );
  NOR4_X1 U373 ( .A1(n1344), .A2(n1345), .A3(n1346), .A4(n1347), .ZN(n1348) );
  NAND4_X1 U374 ( .A1(n1334), .A2(n1339), .A3(n1343), .A4(n1348), .ZN(n1349)
         );
  AOI22_X1 U375 ( .A1(lo_out[10]), .A2(n2281), .B1(n2282), .B2(n1349), .ZN(
        n1350) );
  OAI21_X1 U376 ( .B1(n2283), .B2(n1629), .A(n1350), .ZN(rp1[10]) );
  OAI22_X1 U377 ( .A1(n873), .A2(n3778), .B1(n457), .B2(n3766), .ZN(n1351) );
  OAI22_X1 U378 ( .A1(n393), .A2(n3780), .B1(n361), .B2(n3776), .ZN(n1352) );
  OAI22_X1 U379 ( .A1(n297), .A2(n3764), .B1(n745), .B2(n3768), .ZN(n1353) );
  OAI22_X1 U380 ( .A1(n265), .A2(n3775), .B1(n617), .B2(n3755), .ZN(n1354) );
  NOR4_X1 U381 ( .A1(n1351), .A2(n1352), .A3(n1353), .A4(n1354), .ZN(n1355) );
  OAI22_X1 U382 ( .A1(n809), .A2(n3754), .B1(n329), .B2(n3777), .ZN(n1356) );
  OAI22_X1 U383 ( .A1(n713), .A2(n3762), .B1(n425), .B2(n3760), .ZN(n1357) );
  OAI22_X1 U384 ( .A1(n681), .A2(n3765), .B1(n233), .B2(n3781), .ZN(n1358) );
  OAI22_X1 U385 ( .A1(n9), .A2(n3770), .B1(n585), .B2(n3759), .ZN(n1359) );
  NOR4_X1 U386 ( .A1(n1356), .A2(n1357), .A3(n1358), .A4(n1359), .ZN(n1360) );
  OAI222_X1 U387 ( .A1(n41), .A2(n3773), .B1(n553), .B2(n3782), .C1(n489), 
        .C2(n3757), .ZN(n1361) );
  OAI22_X1 U388 ( .A1(n841), .A2(n3767), .B1(n521), .B2(n3779), .ZN(n1362) );
  OAI22_X1 U389 ( .A1(n777), .A2(n3772), .B1(n649), .B2(n3756), .ZN(n1363) );
  NOR3_X1 U390 ( .A1(n1361), .A2(n1362), .A3(n1363), .ZN(n1364) );
  OAI22_X1 U391 ( .A1(n105), .A2(n3774), .B1(n905), .B2(n3783), .ZN(n1365) );
  OAI22_X1 U392 ( .A1(n137), .A2(n3769), .B1(n937), .B2(n3784), .ZN(n1366) );
  OAI22_X1 U393 ( .A1(n201), .A2(n3758), .B1(n169), .B2(n3761), .ZN(n1367) );
  OAI22_X1 U394 ( .A1(n969), .A2(n3771), .B1(n73), .B2(n3763), .ZN(n1368) );
  NOR4_X1 U395 ( .A1(n1365), .A2(n1366), .A3(n1367), .A4(n1368), .ZN(n1369) );
  NAND4_X1 U396 ( .A1(n1355), .A2(n1360), .A3(n1364), .A4(n1369), .ZN(n1370)
         );
  AOI22_X1 U397 ( .A1(lo_out[8]), .A2(n3786), .B1(n1684), .B2(n1370), .ZN(
        n1371) );
  OAI21_X1 U398 ( .B1(n1626), .B2(n3787), .A(n1371), .ZN(rp2[8]) );
  OAI22_X1 U399 ( .A1(n262), .A2(n2252), .B1(n838), .B2(n2261), .ZN(n1372) );
  OAI22_X1 U400 ( .A1(n102), .A2(n2274), .B1(n6), .B2(n2264), .ZN(n1373) );
  OAI22_X1 U401 ( .A1(n358), .A2(n2260), .B1(n614), .B2(n1678), .ZN(n1374) );
  OAI22_X1 U402 ( .A1(n38), .A2(n2255), .B1(n390), .B2(n2270), .ZN(n1375) );
  NOR4_X1 U403 ( .A1(n1372), .A2(n1373), .A3(n1374), .A4(n1375), .ZN(n1376) );
  OAI22_X1 U404 ( .A1(n646), .A2(n2278), .B1(n678), .B2(n2262), .ZN(n1377) );
  OAI22_X1 U405 ( .A1(n326), .A2(n2256), .B1(n166), .B2(n2257), .ZN(n1378) );
  OAI22_X1 U406 ( .A1(n294), .A2(n2280), .B1(n582), .B2(n2250), .ZN(n1379) );
  OAI22_X1 U407 ( .A1(n870), .A2(n2275), .B1(n486), .B2(n2259), .ZN(n1380) );
  NOR4_X1 U408 ( .A1(n1377), .A2(n1378), .A3(n1379), .A4(n1380), .ZN(n1381) );
  OAI222_X1 U409 ( .A1(n966), .A2(n2258), .B1(n454), .B2(n2268), .C1(n710), 
        .C2(n2269), .ZN(n1382) );
  OAI22_X1 U410 ( .A1(n70), .A2(n2251), .B1(n806), .B2(n2273), .ZN(n1383) );
  OAI22_X1 U411 ( .A1(n422), .A2(n2267), .B1(n230), .B2(n2263), .ZN(n1384) );
  NOR3_X1 U412 ( .A1(n1382), .A2(n1383), .A3(n1384), .ZN(n1385) );
  OAI22_X1 U413 ( .A1(n902), .A2(n2272), .B1(n742), .B2(n2276), .ZN(n1386) );
  OAI22_X1 U414 ( .A1(n198), .A2(n2266), .B1(n518), .B2(n2253), .ZN(n1387) );
  OAI22_X1 U415 ( .A1(n774), .A2(n2279), .B1(n550), .B2(n2265), .ZN(n1388) );
  OAI22_X1 U416 ( .A1(n934), .A2(n2277), .B1(n134), .B2(n1677), .ZN(n1389) );
  NOR4_X1 U417 ( .A1(n1386), .A2(n1387), .A3(n1388), .A4(n1389), .ZN(n1390) );
  NAND4_X1 U418 ( .A1(n1376), .A2(n1381), .A3(n1385), .A4(n1390), .ZN(n1391)
         );
  AOI22_X1 U419 ( .A1(lo_out[5]), .A2(n1679), .B1(n1680), .B2(n1391), .ZN(
        n1392) );
  OAI21_X1 U420 ( .B1(n2283), .B2(n1623), .A(n1392), .ZN(rp1[5]) );
  OAI22_X1 U421 ( .A1(n7), .A2(n3770), .B1(n231), .B2(n3781), .ZN(n1393) );
  OAI22_X1 U422 ( .A1(n359), .A2(n3776), .B1(n711), .B2(n3762), .ZN(n1394) );
  OAI22_X1 U423 ( .A1(n519), .A2(n3779), .B1(n103), .B2(n3774), .ZN(n1395) );
  OAI22_X1 U424 ( .A1(n295), .A2(n3764), .B1(n391), .B2(n1683), .ZN(n1396) );
  NOR4_X1 U425 ( .A1(n1393), .A2(n1394), .A3(n1395), .A4(n1396), .ZN(n1397) );
  OAI22_X1 U426 ( .A1(n167), .A2(n3761), .B1(n871), .B2(n3778), .ZN(n1398) );
  OAI22_X1 U427 ( .A1(n135), .A2(n3769), .B1(n455), .B2(n3766), .ZN(n1399) );
  OAI22_X1 U428 ( .A1(n199), .A2(n3758), .B1(n327), .B2(n3777), .ZN(n1400) );
  OAI22_X1 U429 ( .A1(n775), .A2(n3772), .B1(n743), .B2(n3768), .ZN(n1401) );
  NOR4_X1 U430 ( .A1(n1398), .A2(n1399), .A3(n1400), .A4(n1401), .ZN(n1402) );
  OAI222_X1 U431 ( .A1(n839), .A2(n3767), .B1(n647), .B2(n3756), .C1(n615), 
        .C2(n1681), .ZN(n1403) );
  OAI22_X1 U432 ( .A1(n903), .A2(n3783), .B1(n583), .B2(n3759), .ZN(n1404) );
  OAI22_X1 U433 ( .A1(n487), .A2(n3757), .B1(n71), .B2(n3763), .ZN(n1405) );
  NOR3_X1 U434 ( .A1(n1403), .A2(n1404), .A3(n1405), .ZN(n1406) );
  OAI22_X1 U435 ( .A1(n967), .A2(n3771), .B1(n39), .B2(n3773), .ZN(n1407) );
  OAI22_X1 U436 ( .A1(n263), .A2(n3775), .B1(n679), .B2(n3765), .ZN(n1408) );
  OAI22_X1 U437 ( .A1(n551), .A2(n3782), .B1(n423), .B2(n3760), .ZN(n1409) );
  OAI22_X1 U438 ( .A1(n935), .A2(n3784), .B1(n807), .B2(n3754), .ZN(n1410) );
  NOR4_X1 U439 ( .A1(n1407), .A2(n1408), .A3(n1409), .A4(n1410), .ZN(n1411) );
  NAND4_X1 U440 ( .A1(n1397), .A2(n1402), .A3(n1406), .A4(n1411), .ZN(n1412)
         );
  AOI22_X1 U441 ( .A1(lo_out[6]), .A2(n3786), .B1(n1684), .B2(n1412), .ZN(
        n1413) );
  OAI21_X1 U442 ( .B1(n1624), .B2(n3787), .A(n1413), .ZN(rp2[6]) );
  OAI22_X1 U443 ( .A1(n67), .A2(n2251), .B1(n387), .B2(n2270), .ZN(n1414) );
  OAI22_X1 U444 ( .A1(n195), .A2(n2266), .B1(n227), .B2(n2263), .ZN(n1415) );
  OAI22_X1 U445 ( .A1(n963), .A2(n2258), .B1(n259), .B2(n2252), .ZN(n1416) );
  OAI22_X1 U446 ( .A1(n419), .A2(n2267), .B1(n707), .B2(n2269), .ZN(n1417) );
  NOR4_X1 U447 ( .A1(n1414), .A2(n1415), .A3(n1416), .A4(n1417), .ZN(n1418) );
  OAI22_X1 U448 ( .A1(n3), .A2(n2264), .B1(n451), .B2(n2268), .ZN(n1419) );
  OAI22_X1 U449 ( .A1(n515), .A2(n2253), .B1(n323), .B2(n2256), .ZN(n1420) );
  OAI22_X1 U450 ( .A1(n163), .A2(n2257), .B1(n131), .B2(n2254), .ZN(n1421) );
  OAI22_X1 U451 ( .A1(n835), .A2(n2261), .B1(n771), .B2(n2279), .ZN(n1422) );
  NOR4_X1 U452 ( .A1(n1419), .A2(n1420), .A3(n1421), .A4(n1422), .ZN(n1423) );
  OAI222_X1 U453 ( .A1(n35), .A2(n2255), .B1(n739), .B2(n2276), .C1(n483), 
        .C2(n2259), .ZN(n1424) );
  OAI22_X1 U454 ( .A1(n547), .A2(n2265), .B1(n899), .B2(n2272), .ZN(n1425) );
  OAI22_X1 U455 ( .A1(n99), .A2(n2274), .B1(n291), .B2(n2280), .ZN(n1426) );
  NOR3_X1 U456 ( .A1(n1424), .A2(n1425), .A3(n1426), .ZN(n1427) );
  OAI22_X1 U457 ( .A1(n803), .A2(n2273), .B1(n611), .B2(n2271), .ZN(n1428) );
  OAI22_X1 U458 ( .A1(n931), .A2(n2277), .B1(n867), .B2(n2275), .ZN(n1429) );
  OAI22_X1 U459 ( .A1(n355), .A2(n2260), .B1(n675), .B2(n2262), .ZN(n1430) );
  OAI22_X1 U460 ( .A1(n643), .A2(n2278), .B1(n579), .B2(n2250), .ZN(n1431) );
  NOR4_X1 U461 ( .A1(n1428), .A2(n1429), .A3(n1430), .A4(n1431), .ZN(n1432) );
  NAND4_X1 U462 ( .A1(n1418), .A2(n1423), .A3(n1427), .A4(n1432), .ZN(n1433)
         );
  AOI22_X1 U463 ( .A1(lo_out[2]), .A2(n1679), .B1(n1680), .B2(n1433), .ZN(
        n1434) );
  OAI21_X1 U464 ( .B1(n2283), .B2(n1653), .A(n1434), .ZN(rp1[2]) );
  OAI22_X1 U465 ( .A1(n773), .A2(n3772), .B1(n5), .B2(n3770), .ZN(n1435) );
  OAI22_X1 U466 ( .A1(n741), .A2(n3768), .B1(n677), .B2(n3765), .ZN(n1436) );
  OAI22_X1 U467 ( .A1(n357), .A2(n3776), .B1(n933), .B2(n3784), .ZN(n1437) );
  OAI22_X1 U468 ( .A1(n389), .A2(n1683), .B1(n549), .B2(n3782), .ZN(n1438) );
  NOR4_X1 U469 ( .A1(n1435), .A2(n1436), .A3(n1437), .A4(n1438), .ZN(n1439) );
  OAI22_X1 U470 ( .A1(n261), .A2(n3775), .B1(n197), .B2(n3758), .ZN(n1440) );
  OAI22_X1 U471 ( .A1(n325), .A2(n3777), .B1(n165), .B2(n3761), .ZN(n1441) );
  OAI22_X1 U472 ( .A1(n69), .A2(n3763), .B1(n613), .B2(n3755), .ZN(n1442) );
  OAI22_X1 U473 ( .A1(n517), .A2(n3779), .B1(n133), .B2(n1682), .ZN(n1443) );
  NOR4_X1 U474 ( .A1(n1440), .A2(n1441), .A3(n1442), .A4(n1443), .ZN(n1444) );
  OAI222_X1 U475 ( .A1(n581), .A2(n3759), .B1(n453), .B2(n3766), .C1(n485), 
        .C2(n3757), .ZN(n1445) );
  OAI22_X1 U476 ( .A1(n645), .A2(n3756), .B1(n229), .B2(n3781), .ZN(n1446) );
  OAI22_X1 U477 ( .A1(n293), .A2(n3764), .B1(n709), .B2(n3762), .ZN(n1447) );
  NOR3_X1 U478 ( .A1(n1445), .A2(n1446), .A3(n1447), .ZN(n1448) );
  OAI22_X1 U479 ( .A1(n101), .A2(n3774), .B1(n805), .B2(n3754), .ZN(n1449) );
  OAI22_X1 U480 ( .A1(n965), .A2(n3771), .B1(n421), .B2(n3760), .ZN(n1450) );
  OAI22_X1 U481 ( .A1(n37), .A2(n3773), .B1(n901), .B2(n3783), .ZN(n1451) );
  OAI22_X1 U482 ( .A1(n869), .A2(n3778), .B1(n837), .B2(n3767), .ZN(n1452) );
  NOR4_X1 U483 ( .A1(n1449), .A2(n1450), .A3(n1451), .A4(n1452), .ZN(n1453) );
  NAND4_X1 U484 ( .A1(n1439), .A2(n1444), .A3(n1448), .A4(n1453), .ZN(n1454)
         );
  AOI22_X1 U485 ( .A1(lo_out[4]), .A2(n1685), .B1(n1684), .B2(n1454), .ZN(
        n1455) );
  OAI21_X1 U486 ( .B1(n1649), .B2(n3787), .A(n1455), .ZN(rp2[4]) );
  OAI22_X1 U487 ( .A1(n712), .A2(n2269), .B1(n200), .B2(n2266), .ZN(n1456) );
  OAI22_X1 U488 ( .A1(n744), .A2(n2276), .B1(n616), .B2(n1678), .ZN(n1457) );
  OAI22_X1 U489 ( .A1(n456), .A2(n2268), .B1(n648), .B2(n2278), .ZN(n1458) );
  OAI22_X1 U490 ( .A1(n264), .A2(n2252), .B1(n840), .B2(n2261), .ZN(n1459) );
  NOR4_X1 U491 ( .A1(n1456), .A2(n1457), .A3(n1458), .A4(n1459), .ZN(n1460) );
  OAI22_X1 U492 ( .A1(n488), .A2(n2259), .B1(n392), .B2(n2270), .ZN(n1461) );
  OAI22_X1 U493 ( .A1(n552), .A2(n2265), .B1(n936), .B2(n2277), .ZN(n1462) );
  OAI22_X1 U494 ( .A1(n104), .A2(n2274), .B1(n424), .B2(n2267), .ZN(n1463) );
  OAI22_X1 U495 ( .A1(n520), .A2(n2253), .B1(n776), .B2(n2279), .ZN(n1464) );
  NOR4_X1 U496 ( .A1(n1461), .A2(n1462), .A3(n1463), .A4(n1464), .ZN(n1465) );
  OAI222_X1 U497 ( .A1(n680), .A2(n2262), .B1(n40), .B2(n2255), .C1(n584), 
        .C2(n2250), .ZN(n1466) );
  OAI22_X1 U498 ( .A1(n904), .A2(n2272), .B1(n8), .B2(n2264), .ZN(n1467) );
  OAI22_X1 U499 ( .A1(n168), .A2(n2257), .B1(n328), .B2(n2256), .ZN(n1468) );
  NOR3_X1 U500 ( .A1(n1466), .A2(n1467), .A3(n1468), .ZN(n1469) );
  OAI22_X1 U501 ( .A1(n872), .A2(n2275), .B1(n360), .B2(n2260), .ZN(n1470) );
  OAI22_X1 U502 ( .A1(n72), .A2(n2251), .B1(n968), .B2(n2258), .ZN(n1471) );
  OAI22_X1 U503 ( .A1(n296), .A2(n2280), .B1(n808), .B2(n2273), .ZN(n1472) );
  OAI22_X1 U504 ( .A1(n232), .A2(n2263), .B1(n136), .B2(n1677), .ZN(n1473) );
  NOR4_X1 U505 ( .A1(n1470), .A2(n1471), .A3(n1472), .A4(n1473), .ZN(n1474) );
  NAND4_X1 U506 ( .A1(n1460), .A2(n1465), .A3(n1469), .A4(n1474), .ZN(n1475)
         );
  AOI22_X1 U507 ( .A1(lo_out[7]), .A2(n1679), .B1(n1680), .B2(n1475), .ZN(
        n1476) );
  OAI21_X1 U508 ( .B1(n2283), .B2(n1625), .A(n1476), .ZN(rp1[7]) );
  OAI22_X1 U509 ( .A1(n422), .A2(n3760), .B1(n678), .B2(n3765), .ZN(n1477) );
  OAI22_X1 U510 ( .A1(n6), .A2(n3770), .B1(n966), .B2(n3771), .ZN(n1478) );
  OAI22_X1 U511 ( .A1(n38), .A2(n3773), .B1(n774), .B2(n3772), .ZN(n1479) );
  OAI22_X1 U512 ( .A1(n870), .A2(n3778), .B1(n902), .B2(n3783), .ZN(n1480) );
  NOR4_X1 U513 ( .A1(n1477), .A2(n1478), .A3(n1479), .A4(n1480), .ZN(n1481) );
  OAI22_X1 U514 ( .A1(n550), .A2(n3782), .B1(n70), .B2(n3763), .ZN(n1482) );
  OAI22_X1 U515 ( .A1(n390), .A2(n1683), .B1(n326), .B2(n3777), .ZN(n1483) );
  OAI22_X1 U516 ( .A1(n614), .A2(n1681), .B1(n166), .B2(n3761), .ZN(n1484) );
  OAI22_X1 U517 ( .A1(n486), .A2(n3757), .B1(n102), .B2(n3774), .ZN(n1485) );
  NOR4_X1 U518 ( .A1(n1482), .A2(n1483), .A3(n1484), .A4(n1485), .ZN(n1486) );
  OAI222_X1 U519 ( .A1(n230), .A2(n3781), .B1(n582), .B2(n3759), .C1(n198), 
        .C2(n3758), .ZN(n1487) );
  OAI22_X1 U520 ( .A1(n806), .A2(n3754), .B1(n742), .B2(n3768), .ZN(n1488) );
  OAI22_X1 U521 ( .A1(n710), .A2(n3762), .B1(n262), .B2(n3775), .ZN(n1489) );
  NOR3_X1 U522 ( .A1(n1487), .A2(n1488), .A3(n1489), .ZN(n1490) );
  OAI22_X1 U523 ( .A1(n294), .A2(n3764), .B1(n838), .B2(n3767), .ZN(n1491) );
  OAI22_X1 U524 ( .A1(n934), .A2(n3784), .B1(n358), .B2(n3776), .ZN(n1492) );
  OAI22_X1 U525 ( .A1(n134), .A2(n1682), .B1(n518), .B2(n3779), .ZN(n1493) );
  OAI22_X1 U526 ( .A1(n454), .A2(n3766), .B1(n646), .B2(n3756), .ZN(n1494) );
  NOR4_X1 U527 ( .A1(n1491), .A2(n1492), .A3(n1493), .A4(n1494), .ZN(n1495) );
  NAND4_X1 U528 ( .A1(n1481), .A2(n1486), .A3(n1490), .A4(n1495), .ZN(n1496)
         );
  AOI22_X1 U529 ( .A1(lo_out[5]), .A2(n1685), .B1(n1684), .B2(n1496), .ZN(
        n1497) );
  OAI21_X1 U530 ( .B1(n1623), .B2(n3787), .A(n1497), .ZN(rp2[5]) );
  OAI22_X1 U531 ( .A1(n482), .A2(n2259), .B1(n802), .B2(n2273), .ZN(n1498) );
  OAI22_X1 U532 ( .A1(n418), .A2(n2267), .B1(n130), .B2(n2254), .ZN(n1499) );
  OAI22_X1 U533 ( .A1(n290), .A2(n2280), .B1(n738), .B2(n2276), .ZN(n1500) );
  OAI22_X1 U534 ( .A1(n866), .A2(n2275), .B1(n610), .B2(n2271), .ZN(n1501) );
  NOR4_X1 U535 ( .A1(n1498), .A2(n1499), .A3(n1500), .A4(n1501), .ZN(n1502) );
  OAI22_X1 U536 ( .A1(n450), .A2(n2268), .B1(n546), .B2(n2265), .ZN(n1503) );
  OAI22_X1 U537 ( .A1(n514), .A2(n2253), .B1(n706), .B2(n2269), .ZN(n1504) );
  OAI22_X1 U538 ( .A1(n834), .A2(n2261), .B1(n770), .B2(n2279), .ZN(n1505) );
  OAI22_X1 U539 ( .A1(n66), .A2(n2251), .B1(n2), .B2(n2264), .ZN(n1506) );
  NOR4_X1 U540 ( .A1(n1503), .A2(n1504), .A3(n1505), .A4(n1506), .ZN(n1507) );
  OAI222_X1 U541 ( .A1(n322), .A2(n2256), .B1(n642), .B2(n2278), .C1(n162), 
        .C2(n2257), .ZN(n1508) );
  OAI22_X1 U542 ( .A1(n674), .A2(n2262), .B1(n962), .B2(n2258), .ZN(n1509) );
  OAI22_X1 U543 ( .A1(n578), .A2(n2250), .B1(n98), .B2(n2274), .ZN(n1510) );
  NOR3_X1 U544 ( .A1(n1508), .A2(n1509), .A3(n1510), .ZN(n1511) );
  OAI22_X1 U545 ( .A1(n226), .A2(n2263), .B1(n386), .B2(n2270), .ZN(n1512) );
  OAI22_X1 U546 ( .A1(n34), .A2(n2255), .B1(n354), .B2(n2260), .ZN(n1513) );
  OAI22_X1 U547 ( .A1(n898), .A2(n2272), .B1(n930), .B2(n2277), .ZN(n1514) );
  OAI22_X1 U548 ( .A1(n258), .A2(n2252), .B1(n194), .B2(n2266), .ZN(n1515) );
  NOR4_X1 U549 ( .A1(n1512), .A2(n1513), .A3(n1514), .A4(n1515), .ZN(n1516) );
  NAND4_X1 U550 ( .A1(n1502), .A2(n1507), .A3(n1511), .A4(n1516), .ZN(n1517)
         );
  AOI22_X1 U551 ( .A1(lo_out[1]), .A2(n1679), .B1(n1680), .B2(n1517), .ZN(
        n1518) );
  OAI21_X1 U552 ( .B1(n2283), .B2(n1651), .A(n1518), .ZN(rp1[1]) );
  OAI22_X1 U553 ( .A1(n292), .A2(n3764), .B1(n484), .B2(n3757), .ZN(n1519) );
  OAI22_X1 U554 ( .A1(n772), .A2(n3772), .B1(n420), .B2(n3760), .ZN(n1520) );
  OAI22_X1 U555 ( .A1(n964), .A2(n3771), .B1(n228), .B2(n3781), .ZN(n1521) );
  OAI22_X1 U556 ( .A1(n36), .A2(n3773), .B1(n260), .B2(n3775), .ZN(n1522) );
  NOR4_X1 U557 ( .A1(n1519), .A2(n1520), .A3(n1521), .A4(n1522), .ZN(n1523) );
  OAI22_X1 U558 ( .A1(n196), .A2(n3758), .B1(n708), .B2(n3762), .ZN(n1524) );
  OAI22_X1 U559 ( .A1(n388), .A2(n3780), .B1(n4), .B2(n3770), .ZN(n1525) );
  OAI22_X1 U560 ( .A1(n164), .A2(n3761), .B1(n932), .B2(n3784), .ZN(n1526) );
  OAI22_X1 U561 ( .A1(n740), .A2(n3768), .B1(n676), .B2(n3765), .ZN(n1527) );
  NOR4_X1 U562 ( .A1(n1524), .A2(n1525), .A3(n1526), .A4(n1527), .ZN(n1528) );
  OAI222_X1 U563 ( .A1(n356), .A2(n3776), .B1(n100), .B2(n3774), .C1(n132), 
        .C2(n3769), .ZN(n1529) );
  OAI22_X1 U564 ( .A1(n548), .A2(n3782), .B1(n644), .B2(n3756), .ZN(n1530) );
  OAI22_X1 U565 ( .A1(n612), .A2(n3755), .B1(n68), .B2(n3763), .ZN(n1531) );
  NOR3_X1 U566 ( .A1(n1529), .A2(n1530), .A3(n1531), .ZN(n1532) );
  OAI22_X1 U567 ( .A1(n516), .A2(n3779), .B1(n452), .B2(n3766), .ZN(n1533) );
  OAI22_X1 U568 ( .A1(n324), .A2(n3777), .B1(n804), .B2(n3754), .ZN(n1534) );
  OAI22_X1 U569 ( .A1(n868), .A2(n3778), .B1(n580), .B2(n3759), .ZN(n1535) );
  OAI22_X1 U570 ( .A1(n836), .A2(n3767), .B1(n900), .B2(n3783), .ZN(n1536) );
  NOR4_X1 U571 ( .A1(n1533), .A2(n1534), .A3(n1535), .A4(n1536), .ZN(n1537) );
  NAND4_X1 U572 ( .A1(n1523), .A2(n1528), .A3(n1532), .A4(n1537), .ZN(n1538)
         );
  AOI22_X1 U573 ( .A1(lo_out[3]), .A2(n3786), .B1(n1684), .B2(n1538), .ZN(
        n1539) );
  OAI21_X1 U574 ( .B1(n1648), .B2(n3787), .A(n1539), .ZN(rp2[3]) );
  OAI22_X1 U575 ( .A1(n225), .A2(n2263), .B1(n353), .B2(n2260), .ZN(n1540) );
  OAI22_X1 U576 ( .A1(n641), .A2(n2278), .B1(n161), .B2(n2257), .ZN(n1541) );
  OAI22_X1 U577 ( .A1(n1), .A2(n2264), .B1(n65), .B2(n2251), .ZN(n1542) );
  OAI22_X1 U578 ( .A1(n897), .A2(n2272), .B1(n513), .B2(n2253), .ZN(n1543) );
  NOR4_X1 U579 ( .A1(n1540), .A2(n1541), .A3(n1542), .A4(n1543), .ZN(n1544) );
  OAI22_X1 U580 ( .A1(n545), .A2(n2265), .B1(n97), .B2(n2274), .ZN(n1545) );
  OAI22_X1 U581 ( .A1(n769), .A2(n2279), .B1(n385), .B2(n2270), .ZN(n1546) );
  OAI22_X1 U582 ( .A1(n577), .A2(n2250), .B1(n129), .B2(n1677), .ZN(n1547) );
  OAI22_X1 U583 ( .A1(n33), .A2(n2255), .B1(n417), .B2(n2267), .ZN(n1548) );
  NOR4_X1 U584 ( .A1(n1545), .A2(n1546), .A3(n1547), .A4(n1548), .ZN(n1549) );
  OAI222_X1 U585 ( .A1(n609), .A2(n2271), .B1(n737), .B2(n2276), .C1(n865), 
        .C2(n2275), .ZN(n1550) );
  OAI22_X1 U586 ( .A1(n449), .A2(n2268), .B1(n929), .B2(n2277), .ZN(n1551) );
  OAI22_X1 U587 ( .A1(n321), .A2(n2256), .B1(n833), .B2(n2261), .ZN(n1552) );
  NOR3_X1 U588 ( .A1(n1550), .A2(n1551), .A3(n1552), .ZN(n1553) );
  OAI22_X1 U589 ( .A1(n289), .A2(n2280), .B1(n193), .B2(n2266), .ZN(n1554) );
  OAI22_X1 U590 ( .A1(n481), .A2(n2259), .B1(n961), .B2(n2258), .ZN(n1555) );
  OAI22_X1 U591 ( .A1(n705), .A2(n2269), .B1(n801), .B2(n2273), .ZN(n1556) );
  OAI22_X1 U592 ( .A1(n257), .A2(n2252), .B1(n673), .B2(n2262), .ZN(n1557) );
  NOR4_X1 U593 ( .A1(n1554), .A2(n1555), .A3(n1556), .A4(n1557), .ZN(n1558) );
  NAND4_X1 U594 ( .A1(n1544), .A2(n1549), .A3(n1553), .A4(n1558), .ZN(n1559)
         );
  AOI22_X1 U595 ( .A1(n1679), .A2(lo_out[0]), .B1(n1680), .B2(n1559), .ZN(
        n1560) );
  OAI21_X1 U596 ( .B1(n1628), .B2(n2283), .A(n1560), .ZN(rp1[0]) );
  OAI22_X1 U597 ( .A1(n899), .A2(n3783), .B1(n579), .B2(n3759), .ZN(n1561) );
  OAI22_X1 U598 ( .A1(n291), .A2(n3764), .B1(n803), .B2(n3754), .ZN(n1562) );
  OAI22_X1 U599 ( .A1(n419), .A2(n3760), .B1(n515), .B2(n3779), .ZN(n1563) );
  OAI22_X1 U600 ( .A1(n643), .A2(n3756), .B1(n835), .B2(n3767), .ZN(n1564) );
  NOR4_X1 U601 ( .A1(n1561), .A2(n1562), .A3(n1563), .A4(n1564), .ZN(n1565) );
  OAI22_X1 U602 ( .A1(n259), .A2(n3775), .B1(n771), .B2(n3772), .ZN(n1566) );
  OAI22_X1 U603 ( .A1(n547), .A2(n3782), .B1(n323), .B2(n3777), .ZN(n1567) );
  OAI22_X1 U604 ( .A1(n387), .A2(n1683), .B1(n67), .B2(n3763), .ZN(n1568) );
  OAI22_X1 U605 ( .A1(n99), .A2(n3774), .B1(n931), .B2(n3784), .ZN(n1569) );
  NOR4_X1 U606 ( .A1(n1566), .A2(n1567), .A3(n1568), .A4(n1569), .ZN(n1570) );
  OAI222_X1 U607 ( .A1(n867), .A2(n3778), .B1(n675), .B2(n3765), .C1(n163), 
        .C2(n3761), .ZN(n1571) );
  OAI22_X1 U608 ( .A1(n611), .A2(n3755), .B1(n131), .B2(n1682), .ZN(n1572) );
  OAI22_X1 U609 ( .A1(n707), .A2(n3762), .B1(n451), .B2(n3766), .ZN(n1573) );
  NOR3_X1 U610 ( .A1(n1571), .A2(n1572), .A3(n1573), .ZN(n1574) );
  OAI22_X1 U611 ( .A1(n483), .A2(n3757), .B1(n227), .B2(n3781), .ZN(n1575) );
  OAI22_X1 U612 ( .A1(n355), .A2(n3776), .B1(n195), .B2(n3758), .ZN(n1576) );
  OAI22_X1 U613 ( .A1(n739), .A2(n3768), .B1(n35), .B2(n3773), .ZN(n1577) );
  OAI22_X1 U614 ( .A1(n963), .A2(n3771), .B1(n3), .B2(n3770), .ZN(n1578) );
  NOR4_X1 U615 ( .A1(n1575), .A2(n1576), .A3(n1577), .A4(n1578), .ZN(n1579) );
  NAND4_X1 U616 ( .A1(n1565), .A2(n1570), .A3(n1574), .A4(n1579), .ZN(n1580)
         );
  AOI22_X1 U617 ( .A1(lo_out[2]), .A2(n3786), .B1(n3785), .B2(n1580), .ZN(
        n1581) );
  OAI21_X1 U618 ( .B1(n1653), .B2(n3787), .A(n1581), .ZN(rp2[2]) );
  INV_X2 U619 ( .A(hilo_wr_en), .ZN(n1688) );
  BUF_X1 U620 ( .A(n1688), .Z(n1582) );
  BUF_X1 U621 ( .A(n1688), .Z(n1615) );
  BUF_X1 U622 ( .A(n1710), .Z(n1588) );
  BUF_X1 U623 ( .A(n1696), .Z(n1587) );
  BUF_X1 U624 ( .A(n1782), .Z(n1584) );
  BUF_X1 U625 ( .A(n1738), .Z(n1583) );
  BUF_X1 U626 ( .A(n1692), .Z(n1589) );
  BUF_X1 U627 ( .A(n1764), .Z(n1591) );
  BUF_X1 U628 ( .A(n1798), .Z(n1586) );
  BUF_X1 U629 ( .A(n1726), .Z(n1590) );
  BUF_X1 U630 ( .A(n1752), .Z(n1585) );
  BUF_X1 U631 ( .A(n1702), .Z(n1593) );
  BUF_X1 U632 ( .A(n1732), .Z(n1611) );
  BUF_X1 U633 ( .A(n1790), .Z(n1601) );
  BUF_X1 U634 ( .A(n1755), .Z(n1607) );
  BUF_X1 U635 ( .A(n1742), .Z(n1603) );
  BUF_X1 U636 ( .A(n1794), .Z(n1596) );
  BUF_X1 U637 ( .A(n1786), .Z(n1606) );
  BUF_X1 U638 ( .A(n1758), .Z(n1608) );
  BUF_X1 U639 ( .A(n1778), .Z(n1609) );
  BUF_X1 U640 ( .A(n1746), .Z(n1602) );
  BUF_X1 U641 ( .A(n1699), .Z(n1594) );
  BUF_X1 U642 ( .A(n1693), .Z(n1600) );
  BUF_X1 U643 ( .A(n1716), .Z(n1595) );
  BUF_X1 U644 ( .A(n1768), .Z(n1605) );
  BUF_X1 U645 ( .A(n1774), .Z(n1612) );
  BUF_X1 U646 ( .A(n1729), .Z(n1597) );
  BUF_X1 U647 ( .A(n1706), .Z(n1599) );
  BUF_X1 U648 ( .A(n1735), .Z(n1604) );
  BUF_X1 U649 ( .A(n1749), .Z(n1610) );
  BUF_X1 U650 ( .A(n1761), .Z(n1613) );
  BUF_X1 U651 ( .A(n1835), .Z(n1592) );
  BUF_X1 U652 ( .A(n1723), .Z(n1598) );
  BUF_X1 U653 ( .A(n1720), .Z(n1614) );
  INV_X2 U654 ( .A(wp[0]), .ZN(n1802) );
  INV_X2 U655 ( .A(wp[1]), .ZN(n1803) );
  INV_X2 U656 ( .A(wp[2]), .ZN(n1804) );
  INV_X2 U657 ( .A(wp[3]), .ZN(n1805) );
  INV_X2 U658 ( .A(wp[4]), .ZN(n1806) );
  INV_X2 U659 ( .A(wp[5]), .ZN(n1807) );
  INV_X2 U660 ( .A(wp[6]), .ZN(n1808) );
  INV_X2 U661 ( .A(wp[7]), .ZN(n1809) );
  INV_X2 U662 ( .A(wp[8]), .ZN(n1810) );
  INV_X2 U663 ( .A(wp[9]), .ZN(n1811) );
  INV_X2 U664 ( .A(wp[10]), .ZN(n1812) );
  INV_X2 U665 ( .A(wp[11]), .ZN(n1813) );
  INV_X2 U666 ( .A(wp[12]), .ZN(n1814) );
  INV_X2 U667 ( .A(wp[13]), .ZN(n1815) );
  INV_X2 U668 ( .A(wp[14]), .ZN(n1816) );
  INV_X2 U669 ( .A(wp[15]), .ZN(n1817) );
  INV_X2 U670 ( .A(wp[16]), .ZN(n1818) );
  INV_X2 U671 ( .A(wp[17]), .ZN(n1819) );
  INV_X2 U672 ( .A(wp[18]), .ZN(n1820) );
  INV_X2 U673 ( .A(wp[19]), .ZN(n1821) );
  INV_X2 U674 ( .A(wp[20]), .ZN(n1822) );
  INV_X2 U675 ( .A(wp[21]), .ZN(n1823) );
  INV_X2 U676 ( .A(wp[22]), .ZN(n1824) );
  INV_X2 U677 ( .A(wp[23]), .ZN(n1825) );
  INV_X2 U678 ( .A(wp[24]), .ZN(n1826) );
  INV_X2 U679 ( .A(wp[25]), .ZN(n1827) );
  INV_X2 U680 ( .A(wp[26]), .ZN(n1828) );
  INV_X2 U681 ( .A(wp[27]), .ZN(n1829) );
  BUF_X2 U682 ( .A(n1781), .Z(n1617) );
  BUF_X2 U683 ( .A(n1751), .Z(n1619) );
  BUF_X2 U684 ( .A(n1797), .Z(n1616) );
  BUF_X2 U685 ( .A(n1763), .Z(n1618) );
  BUF_X2 U686 ( .A(n1834), .Z(n1620) );
  BUF_X2 U687 ( .A(n1785), .Z(n1621) );
  NOR3_X1 U688 ( .A1(wp_addr[2]), .A2(wp_addr[1]), .A3(n1703), .ZN(n1776) );
  NAND2_X2 U689 ( .A1(rp1_out_sel[1]), .A2(n1853), .ZN(n2283) );
  BUF_X1 U690 ( .A(n1688), .Z(n1622) );
  NAND2_X2 U691 ( .A1(rp2_out_sel[1]), .A2(n2284), .ZN(n3787) );
  INV_X8 U692 ( .A(clk), .ZN(n993) );
  BUF_X1 U693 ( .A(n1695), .Z(n1655) );
  BUF_X1 U694 ( .A(n1725), .Z(n1662) );
  NAND2_X1 U695 ( .A1(rst), .A2(n1724), .ZN(n1726) );
  NAND2_X1 U696 ( .A1(rst), .A2(n1795), .ZN(n1798) );
  BUF_X1 U697 ( .A(n1737), .Z(n1666) );
  NAND2_X1 U698 ( .A1(rst), .A2(n1750), .ZN(n1752) );
  BUF_X1 U699 ( .A(n1709), .Z(n1659) );
  NAND2_X1 U700 ( .A1(rst), .A2(n1708), .ZN(n1710) );
  NAND2_X1 U701 ( .A1(rst), .A2(n1691), .ZN(n1692) );
  NAND2_X1 U702 ( .A1(rst), .A2(n1762), .ZN(n1764) );
  NAND2_X1 U703 ( .A1(rst), .A2(n1736), .ZN(n1738) );
  NAND2_X1 U704 ( .A1(rst), .A2(n1694), .ZN(n1696) );
  NAND2_X1 U705 ( .A1(rst), .A2(n1779), .ZN(n1782) );
  NAND3_X1 U706 ( .A1(rst), .A2(n1714), .A3(n1780), .ZN(n1695) );
  BUF_X1 U707 ( .A(n1789), .Z(n1675) );
  NAND2_X1 U708 ( .A1(rst), .A2(n1771), .ZN(n1774) );
  NAND2_X1 U709 ( .A1(rst), .A2(n1700), .ZN(n1702) );
  BUF_X1 U710 ( .A(n1728), .Z(n1663) );
  BUF_X1 U711 ( .A(n1741), .Z(n1667) );
  NAND2_X1 U712 ( .A1(rst), .A2(n1721), .ZN(n1723) );
  NAND2_X1 U713 ( .A1(rst), .A2(n1730), .ZN(n1732) );
  NAND2_X1 U714 ( .A1(rst), .A2(n1727), .ZN(n1729) );
  NAND2_X1 U715 ( .A1(rst), .A2(n1739), .ZN(n1742) );
  NAND2_X1 U716 ( .A1(rst), .A2(n1697), .ZN(n1699) );
  NAND2_X1 U717 ( .A1(rst), .A2(n1787), .ZN(n1790) );
  NAND3_X1 U718 ( .A1(rst), .A2(n1780), .A3(n1740), .ZN(n1725) );
  BUF_X1 U719 ( .A(n1754), .Z(n1669) );
  NAND2_X1 U720 ( .A1(rst), .A2(n1791), .ZN(n1794) );
  BUF_X1 U721 ( .A(n1722), .Z(n1661) );
  NAND2_X1 U722 ( .A1(rst), .A2(n1756), .ZN(n1758) );
  NAND2_X1 U723 ( .A1(rst), .A2(n1799), .ZN(n1835) );
  INV_X2 U724 ( .A(wp[30]), .ZN(n1832) );
  NAND2_X1 U725 ( .A1(rst), .A2(n1733), .ZN(n1735) );
  INV_X2 U726 ( .A(wp[29]), .ZN(n1831) );
  BUF_X1 U727 ( .A(n1793), .Z(n1676) );
  INV_X2 U728 ( .A(wp[28]), .ZN(n1830) );
  BUF_X1 U729 ( .A(n1698), .Z(n1656) );
  BUF_X1 U730 ( .A(n1731), .Z(n1664) );
  BUF_X1 U731 ( .A(n1773), .Z(n1673) );
  NAND2_X1 U732 ( .A1(rst), .A2(n1747), .ZN(n1749) );
  BUF_X1 U733 ( .A(n1748), .Z(n1668) );
  INV_X2 U734 ( .A(wp[31]), .ZN(n1833) );
  BUF_X1 U735 ( .A(n1757), .Z(n1670) );
  BUF_X1 U736 ( .A(n1760), .Z(n1671) );
  BUF_X1 U737 ( .A(n1734), .Z(n1665) );
  BUF_X1 U738 ( .A(n1767), .Z(n1672) );
  BUF_X1 U739 ( .A(n1777), .Z(n1674) );
  NAND2_X2 U740 ( .A1(rst), .A2(n1718), .ZN(n1719) );
  NAND2_X1 U741 ( .A1(rst), .A2(n1775), .ZN(n1778) );
  NAND2_X1 U742 ( .A1(rst), .A2(n1783), .ZN(n1786) );
  NAND3_X1 U743 ( .A1(rst), .A2(n1796), .A3(n1740), .ZN(n1737) );
  NAND2_X1 U744 ( .A1(rst), .A2(n1690), .ZN(n1693) );
  NAND2_X1 U745 ( .A1(rst), .A2(n1753), .ZN(n1755) );
  BUF_X1 U746 ( .A(n1715), .Z(n1660) );
  NAND2_X1 U747 ( .A1(rst), .A2(n1765), .ZN(n1768) );
  NAND2_X1 U748 ( .A1(rst), .A2(n1744), .ZN(n1746) );
  NAND2_X1 U749 ( .A1(rst), .A2(n1759), .ZN(n1761) );
  NAND3_X1 U750 ( .A1(rst), .A2(n1714), .A3(n1796), .ZN(n1709) );
  BUF_X1 U751 ( .A(n1701), .Z(n1657) );
  BUF_X1 U752 ( .A(n1705), .Z(n1658) );
  NAND2_X1 U753 ( .A1(rst), .A2(n1704), .ZN(n1706) );
  NAND2_X1 U754 ( .A1(rst), .A2(n1713), .ZN(n1716) );
  NAND3_X1 U755 ( .A1(rst), .A2(n1772), .A3(n1800), .ZN(n1773) );
  NAND3_X1 U756 ( .A1(rst), .A2(n1788), .A3(n1740), .ZN(n1731) );
  NAND3_X1 U757 ( .A1(rst), .A2(n1792), .A3(n1766), .ZN(n1760) );
  NAND3_X1 U758 ( .A1(rst), .A2(n1801), .A3(n1766), .ZN(n1767) );
  NOR2_X1 U759 ( .A1(wp_addr[2]), .A2(n1707), .ZN(n1780) );
  NAND3_X1 U760 ( .A1(rst), .A2(n1776), .A3(n1766), .ZN(n1748) );
  NAND3_X1 U761 ( .A1(rst), .A2(n1788), .A3(n1800), .ZN(n1789) );
  NAND3_X1 U762 ( .A1(rst), .A2(n1792), .A3(n1740), .ZN(n1734) );
  NAND3_X1 U763 ( .A1(rst), .A2(n1776), .A3(n1800), .ZN(n1777) );
  NAND3_X1 U764 ( .A1(rst), .A2(n1792), .A3(n1800), .ZN(n1793) );
  NAND3_X1 U765 ( .A1(rst), .A2(n1714), .A3(n1784), .ZN(n1698) );
  NAND3_X1 U766 ( .A1(rst), .A2(n1788), .A3(n1766), .ZN(n1757) );
  NAND3_X1 U767 ( .A1(rst), .A2(n1714), .A3(n1801), .ZN(n1715) );
  NAND3_X1 U768 ( .A1(rst), .A2(n1784), .A3(n1766), .ZN(n1754) );
  NOR2_X1 U769 ( .A1(n1712), .A2(n1707), .ZN(n1796) );
  NAND3_X1 U770 ( .A1(rst), .A2(n1714), .A3(n1792), .ZN(n1705) );
  NAND2_X1 U771 ( .A1(rst), .A2(n1717), .ZN(n1720) );
  NAND3_X1 U772 ( .A1(rst), .A2(n1801), .A3(n1740), .ZN(n1741) );
  NAND3_X1 U773 ( .A1(rst), .A2(n1776), .A3(n1740), .ZN(n1722) );
  NAND3_X1 U774 ( .A1(rst), .A2(n1784), .A3(n1740), .ZN(n1728) );
  NAND3_X1 U775 ( .A1(rst), .A2(n1714), .A3(n1788), .ZN(n1701) );
  NAND2_X2 U776 ( .A1(n1839), .A2(n1850), .ZN(n2273) );
  NOR2_X1 U777 ( .A1(wp_addr[2]), .A2(n1711), .ZN(n1784) );
  NAND2_X2 U778 ( .A1(n2299), .A2(n2312), .ZN(n3759) );
  NOR2_X2 U779 ( .A1(wp_addr[4]), .A2(n1743), .ZN(n1714) );
  NAND2_X2 U780 ( .A1(n1850), .A2(n1849), .ZN(n2255) );
  NAND2_X2 U781 ( .A1(n1852), .A2(n1843), .ZN(n2268) );
  NAND2_X2 U782 ( .A1(n1850), .A2(n1848), .ZN(n2250) );
  NAND2_X2 U783 ( .A1(n2311), .A2(n2304), .ZN(n3770) );
  NAND2_X2 U784 ( .A1(n1839), .A2(n1852), .ZN(n2277) );
  NAND2_X2 U785 ( .A1(n2307), .A2(n2308), .ZN(n3771) );
  NAND2_X2 U786 ( .A1(n2307), .A2(n2304), .ZN(n3758) );
  NAND2_X2 U787 ( .A1(n2311), .A2(n2306), .ZN(n3757) );
  NAND2_X2 U788 ( .A1(n2298), .A2(n2311), .ZN(n3781) );
  NAND2_X2 U789 ( .A1(n1843), .A2(n1850), .ZN(n2256) );
  NAND2_X2 U790 ( .A1(n1852), .A2(n1844), .ZN(n2258) );
  NAND2_X2 U791 ( .A1(n2307), .A2(n2299), .ZN(n3762) );
  NAND2_X2 U792 ( .A1(n2307), .A2(n2313), .ZN(n3766) );
  NOR2_X2 U793 ( .A1(n1770), .A2(n1769), .ZN(n1800) );
  NAND2_X2 U794 ( .A1(n1842), .A2(n1845), .ZN(n2259) );
  NAND2_X2 U795 ( .A1(n2307), .A2(n2305), .ZN(n3784) );
  NAND2_X2 U796 ( .A1(n2305), .A2(n2310), .ZN(n3778) );
  NAND2_X2 U797 ( .A1(n2307), .A2(n2306), .ZN(n3765) );
  NAND2_X2 U798 ( .A1(n2298), .A2(n2310), .ZN(n3776) );
  NOR2_X1 U799 ( .A1(n1712), .A2(n1711), .ZN(n1801) );
  BUF_X1 U800 ( .A(n2281), .Z(n1679) );
  NAND2_X2 U801 ( .A1(n2310), .A2(n2309), .ZN(n3774) );
  NAND2_X2 U802 ( .A1(n1850), .A2(n1844), .ZN(n2261) );
  NAND2_X2 U803 ( .A1(n1852), .A2(n1851), .ZN(n2267) );
  NAND2_X2 U804 ( .A1(n1852), .A2(n1846), .ZN(n2266) );
  NAND2_X2 U805 ( .A1(n2311), .A2(n2305), .ZN(n3768) );
  NAND2_X2 U806 ( .A1(n1845), .A2(n1848), .ZN(n2253) );
  NAND2_X2 U807 ( .A1(n2311), .A2(n2299), .ZN(n3779) );
  NAND2_X2 U808 ( .A1(n1847), .A2(n1839), .ZN(n2275) );
  NAND2_X2 U809 ( .A1(n1842), .A2(n1852), .ZN(n2262) );
  NAND2_X2 U810 ( .A1(n1850), .A2(n1846), .ZN(n2251) );
  NAND2_X2 U811 ( .A1(n2307), .A2(n2298), .ZN(n3760) );
  NAND2_X2 U812 ( .A1(n2311), .A2(n2308), .ZN(n3772) );
  NAND2_X2 U813 ( .A1(n1845), .A2(n1846), .ZN(n2264) );
  NAND2_X2 U814 ( .A1(n1845), .A2(n1843), .ZN(n2252) );
  NAND2_X2 U815 ( .A1(n1847), .A2(n1848), .ZN(n2278) );
  NAND2_X2 U816 ( .A1(n1845), .A2(n1851), .ZN(n2263) );
  NAND2_X2 U817 ( .A1(n1847), .A2(n1851), .ZN(n2260) );
  NAND2_X2 U818 ( .A1(n2299), .A2(n2310), .ZN(n3756) );
  NAND2_X2 U819 ( .A1(n1845), .A2(n1844), .ZN(n2279) );
  NOR2_X2 U820 ( .A1(n1770), .A2(n1743), .ZN(n1766) );
  NAND2_X2 U821 ( .A1(n1850), .A2(n1851), .ZN(n2280) );
  NAND2_X2 U822 ( .A1(n2310), .A2(n2308), .ZN(n3783) );
  NAND2_X2 U823 ( .A1(n1847), .A2(n1843), .ZN(n2270) );
  NAND2_X2 U824 ( .A1(n1847), .A2(n1849), .ZN(n2274) );
  NAND2_X2 U825 ( .A1(n1842), .A2(n1850), .ZN(n2265) );
  NAND2_X2 U826 ( .A1(n1852), .A2(n1848), .ZN(n2269) );
  NAND2_X2 U827 ( .A1(n1845), .A2(n1839), .ZN(n2276) );
  BUF_X1 U828 ( .A(n3786), .Z(n1685) );
  NAND2_X2 U829 ( .A1(n2311), .A2(n2313), .ZN(n3775) );
  NAND2_X2 U830 ( .A1(n2305), .A2(n2312), .ZN(n3754) );
  NAND2_X2 U831 ( .A1(n1847), .A2(n1844), .ZN(n2272) );
  NAND2_X2 U832 ( .A1(n1852), .A2(n1849), .ZN(n2257) );
  INV_X1 U833 ( .A(n1688), .ZN(n1686) );
  INV_X1 U834 ( .A(n1688), .ZN(n1687) );
  BUF_X1 U835 ( .A(n2282), .Z(n1680) );
  NAND2_X1 U836 ( .A1(wp_en), .A2(n1689), .ZN(n1743) );
  NAND2_X2 U837 ( .A1(n2307), .A2(n2309), .ZN(n3761) );
  NOR3_X2 U838 ( .A1(wp_addr[1]), .A2(n1712), .A3(n1703), .ZN(n1792) );
  NOR3_X2 U839 ( .A1(wp_addr[1]), .A2(wp_addr[0]), .A3(n1712), .ZN(n1788) );
  INV_X1 U840 ( .A(wp_addr[2]), .ZN(n1712) );
  NAND2_X2 U841 ( .A1(n2304), .A2(n2312), .ZN(n3763) );
  NAND2_X2 U842 ( .A1(n2312), .A2(n2308), .ZN(n3767) );
  NAND2_X2 U843 ( .A1(n2306), .A2(n2312), .ZN(n3782) );
  NAND2_X2 U844 ( .A1(n2298), .A2(n2312), .ZN(n3764) );
  NAND2_X2 U845 ( .A1(n2312), .A2(n2309), .ZN(n3773) );
  BUF_X1 U846 ( .A(n3785), .Z(n1684) );
  NAND2_X2 U847 ( .A1(n2313), .A2(n2312), .ZN(n3777) );
  NAND2_X1 U848 ( .A1(wp_addr[1]), .A2(n1703), .ZN(n1707) );
  INV_X1 U849 ( .A(wp_addr[3]), .ZN(n1689) );
  NAND2_X1 U850 ( .A1(wp_en), .A2(wp_addr[3]), .ZN(n1769) );
  INV_X1 U851 ( .A(wp_addr[0]), .ZN(n1703) );
  NOR2_X2 U852 ( .A1(wp_addr[4]), .A2(n1769), .ZN(n1740) );
  INV_X1 U853 ( .A(wp_addr[4]), .ZN(n1770) );
  INV_X1 U854 ( .A(n1717), .ZN(n1718) );
  NOR3_X1 U855 ( .A1(wp_addr[2]), .A2(wp_addr[1]), .A3(wp_addr[0]), .ZN(n1772)
         );
  NAND3_X2 U856 ( .A1(rst), .A2(n1772), .A3(n1766), .ZN(n1745) );
  NAND2_X1 U857 ( .A1(wp_addr[1]), .A2(wp_addr[0]), .ZN(n1711) );
  INV_X1 U858 ( .A(rp2_out_sel[0]), .ZN(n2284) );
  BUF_X1 U859 ( .A(n3769), .Z(n1682) );
  BUF_X1 U860 ( .A(n3780), .Z(n1683) );
  BUF_X1 U861 ( .A(n3755), .Z(n1681) );
  BUF_X1 U862 ( .A(n2271), .Z(n1678) );
  BUF_X1 U863 ( .A(n2254), .Z(n1677) );
  NAND2_X1 U864 ( .A1(n1776), .A2(n1714), .ZN(n1690) );
  INV_X1 U865 ( .A(n1690), .ZN(n1691) );
  OAI22_X1 U866 ( .A1(n1), .A2(n1600), .B1(n1589), .B2(n1802), .ZN(n3614) );
  OAI22_X1 U867 ( .A1(n2), .A2(n1600), .B1(n1803), .B2(n1589), .ZN(n3613) );
  OAI22_X1 U868 ( .A1(n3), .A2(n1600), .B1(n1804), .B2(n1589), .ZN(n3612) );
  OAI22_X1 U869 ( .A1(n4), .A2(n1600), .B1(n1805), .B2(n1589), .ZN(n3611) );
  OAI22_X1 U870 ( .A1(n5), .A2(n1600), .B1(n1806), .B2(n1589), .ZN(n3610) );
  OAI22_X1 U871 ( .A1(n6), .A2(n1600), .B1(n1807), .B2(n1589), .ZN(n3609) );
  OAI22_X1 U872 ( .A1(n7), .A2(n1600), .B1(n1808), .B2(n1589), .ZN(n3608) );
  OAI22_X1 U873 ( .A1(n8), .A2(n1600), .B1(n1809), .B2(n1589), .ZN(n3607) );
  OAI22_X1 U874 ( .A1(n9), .A2(n1600), .B1(n1810), .B2(n1589), .ZN(n3606) );
  OAI22_X1 U875 ( .A1(n10), .A2(n1600), .B1(n1811), .B2(n1589), .ZN(n3605) );
  OAI22_X1 U876 ( .A1(n11), .A2(n1600), .B1(n1812), .B2(n1589), .ZN(n3604) );
  OAI22_X1 U877 ( .A1(n12), .A2(n1600), .B1(n1813), .B2(n1589), .ZN(n3603) );
  OAI22_X1 U878 ( .A1(n13), .A2(n1600), .B1(n1814), .B2(n1589), .ZN(n3602) );
  OAI22_X1 U879 ( .A1(n14), .A2(n1600), .B1(n1815), .B2(n1589), .ZN(n3601) );
  OAI22_X1 U880 ( .A1(n15), .A2(n1600), .B1(n1816), .B2(n1589), .ZN(n3600) );
  OAI22_X1 U881 ( .A1(n16), .A2(n1600), .B1(n1817), .B2(n1589), .ZN(n3599) );
  OAI22_X1 U882 ( .A1(n17), .A2(n1600), .B1(n1818), .B2(n1589), .ZN(n3598) );
  OAI22_X1 U883 ( .A1(n18), .A2(n1600), .B1(n1819), .B2(n1589), .ZN(n3597) );
  OAI22_X1 U884 ( .A1(n19), .A2(n1600), .B1(n1820), .B2(n1589), .ZN(n3596) );
  OAI22_X1 U885 ( .A1(n20), .A2(n1600), .B1(n1821), .B2(n1589), .ZN(n3595) );
  OAI22_X1 U886 ( .A1(n21), .A2(n1600), .B1(n1822), .B2(n1589), .ZN(n3594) );
  OAI22_X1 U887 ( .A1(n22), .A2(n1600), .B1(n1823), .B2(n1589), .ZN(n3593) );
  OAI22_X1 U888 ( .A1(n23), .A2(n1600), .B1(n1824), .B2(n1589), .ZN(n3592) );
  OAI22_X1 U889 ( .A1(n24), .A2(n1600), .B1(n1825), .B2(n1589), .ZN(n3591) );
  OAI22_X1 U890 ( .A1(n25), .A2(n1693), .B1(n1826), .B2(n1692), .ZN(n3590) );
  OAI22_X1 U891 ( .A1(n26), .A2(n1693), .B1(n1827), .B2(n1692), .ZN(n3589) );
  OAI22_X1 U892 ( .A1(n27), .A2(n1693), .B1(n1828), .B2(n1589), .ZN(n3588) );
  OAI22_X1 U893 ( .A1(n28), .A2(n1693), .B1(n1829), .B2(n1589), .ZN(n3587) );
  OAI22_X1 U894 ( .A1(n29), .A2(n1693), .B1(n1830), .B2(n1692), .ZN(n3586) );
  OAI22_X1 U895 ( .A1(n30), .A2(n1693), .B1(n1831), .B2(n1692), .ZN(n3585) );
  OAI22_X1 U896 ( .A1(n31), .A2(n1600), .B1(n1832), .B2(n1692), .ZN(n3584) );
  OAI22_X1 U897 ( .A1(n32), .A2(n1600), .B1(n1833), .B2(n1692), .ZN(n3583) );
  NAND2_X1 U898 ( .A1(n1714), .A2(n1780), .ZN(n1694) );
  OAI22_X1 U899 ( .A1(n33), .A2(n1587), .B1(n1695), .B2(n1802), .ZN(n3582) );
  OAI22_X1 U900 ( .A1(n34), .A2(n1587), .B1(n1695), .B2(n1803), .ZN(n3581) );
  OAI22_X1 U901 ( .A1(n35), .A2(n1587), .B1(n1695), .B2(n1804), .ZN(n3580) );
  OAI22_X1 U902 ( .A1(n36), .A2(n1587), .B1(n1695), .B2(n1805), .ZN(n3579) );
  OAI22_X1 U903 ( .A1(n37), .A2(n1587), .B1(n1695), .B2(n1806), .ZN(n3578) );
  OAI22_X1 U904 ( .A1(n38), .A2(n1587), .B1(n1695), .B2(n1807), .ZN(n3577) );
  OAI22_X1 U905 ( .A1(n39), .A2(n1587), .B1(n1695), .B2(n1808), .ZN(n3576) );
  OAI22_X1 U906 ( .A1(n40), .A2(n1587), .B1(n1695), .B2(n1809), .ZN(n3575) );
  OAI22_X1 U907 ( .A1(n41), .A2(n1587), .B1(n1695), .B2(n1810), .ZN(n3574) );
  OAI22_X1 U908 ( .A1(n42), .A2(n1587), .B1(n1695), .B2(n1811), .ZN(n3573) );
  OAI22_X1 U909 ( .A1(n43), .A2(n1587), .B1(n1695), .B2(n1812), .ZN(n3572) );
  OAI22_X1 U910 ( .A1(n44), .A2(n1587), .B1(n1695), .B2(n1813), .ZN(n3571) );
  OAI22_X1 U911 ( .A1(n45), .A2(n1587), .B1(n1655), .B2(n1814), .ZN(n3570) );
  OAI22_X1 U912 ( .A1(n46), .A2(n1587), .B1(n1655), .B2(n1815), .ZN(n3569) );
  OAI22_X1 U913 ( .A1(n47), .A2(n1587), .B1(n1655), .B2(n1816), .ZN(n3568) );
  OAI22_X1 U914 ( .A1(n48), .A2(n1587), .B1(n1655), .B2(n1817), .ZN(n3567) );
  OAI22_X1 U915 ( .A1(n49), .A2(n1587), .B1(n1655), .B2(n1818), .ZN(n3566) );
  OAI22_X1 U916 ( .A1(n50), .A2(n1587), .B1(n1655), .B2(n1819), .ZN(n3565) );
  OAI22_X1 U917 ( .A1(n51), .A2(n1587), .B1(n1655), .B2(n1820), .ZN(n3564) );
  OAI22_X1 U918 ( .A1(n52), .A2(n1587), .B1(n1655), .B2(n1821), .ZN(n3563) );
  OAI22_X1 U919 ( .A1(n53), .A2(n1587), .B1(n1655), .B2(n1822), .ZN(n3562) );
  OAI22_X1 U920 ( .A1(n54), .A2(n1587), .B1(n1655), .B2(n1823), .ZN(n3561) );
  OAI22_X1 U921 ( .A1(n55), .A2(n1587), .B1(n1655), .B2(n1824), .ZN(n3560) );
  OAI22_X1 U922 ( .A1(n56), .A2(n1587), .B1(n1655), .B2(n1825), .ZN(n3559) );
  OAI22_X1 U923 ( .A1(n57), .A2(n1696), .B1(n1695), .B2(n1826), .ZN(n3558) );
  OAI22_X1 U924 ( .A1(n58), .A2(n1696), .B1(n1655), .B2(n1827), .ZN(n3557) );
  OAI22_X1 U925 ( .A1(n59), .A2(n1696), .B1(n1655), .B2(n1828), .ZN(n3556) );
  OAI22_X1 U926 ( .A1(n60), .A2(n1696), .B1(n1655), .B2(n1829), .ZN(n3555) );
  OAI22_X1 U927 ( .A1(n61), .A2(n1696), .B1(n1695), .B2(n1830), .ZN(n3554) );
  OAI22_X1 U928 ( .A1(n62), .A2(n1696), .B1(n1695), .B2(n1831), .ZN(n3553) );
  OAI22_X1 U929 ( .A1(n63), .A2(n1587), .B1(n1655), .B2(n1832), .ZN(n3552) );
  OAI22_X1 U930 ( .A1(n64), .A2(n1587), .B1(n1655), .B2(n1833), .ZN(n3551) );
  NAND2_X1 U931 ( .A1(n1714), .A2(n1784), .ZN(n1697) );
  OAI22_X1 U932 ( .A1(n65), .A2(n1594), .B1(n1698), .B2(n1802), .ZN(n3550) );
  OAI22_X1 U933 ( .A1(n66), .A2(n1594), .B1(n1698), .B2(n1803), .ZN(n3549) );
  OAI22_X1 U934 ( .A1(n67), .A2(n1594), .B1(n1698), .B2(n1804), .ZN(n3548) );
  OAI22_X1 U935 ( .A1(n68), .A2(n1594), .B1(n1698), .B2(n1805), .ZN(n3547) );
  OAI22_X1 U936 ( .A1(n69), .A2(n1594), .B1(n1698), .B2(n1806), .ZN(n3546) );
  OAI22_X1 U937 ( .A1(n70), .A2(n1594), .B1(n1698), .B2(n1807), .ZN(n3545) );
  OAI22_X1 U938 ( .A1(n71), .A2(n1594), .B1(n1698), .B2(n1808), .ZN(n3544) );
  OAI22_X1 U939 ( .A1(n72), .A2(n1594), .B1(n1698), .B2(n1809), .ZN(n3543) );
  OAI22_X1 U940 ( .A1(n73), .A2(n1594), .B1(n1698), .B2(n1810), .ZN(n3542) );
  OAI22_X1 U941 ( .A1(n74), .A2(n1594), .B1(n1698), .B2(n1811), .ZN(n3541) );
  OAI22_X1 U942 ( .A1(n75), .A2(n1594), .B1(n1698), .B2(n1812), .ZN(n3540) );
  OAI22_X1 U943 ( .A1(n76), .A2(n1594), .B1(n1698), .B2(n1813), .ZN(n3539) );
  OAI22_X1 U944 ( .A1(n77), .A2(n1594), .B1(n1656), .B2(n1814), .ZN(n3538) );
  OAI22_X1 U945 ( .A1(n78), .A2(n1594), .B1(n1656), .B2(n1815), .ZN(n3537) );
  OAI22_X1 U946 ( .A1(n79), .A2(n1594), .B1(n1656), .B2(n1816), .ZN(n3536) );
  OAI22_X1 U947 ( .A1(n80), .A2(n1594), .B1(n1656), .B2(n1817), .ZN(n3535) );
  OAI22_X1 U948 ( .A1(n81), .A2(n1594), .B1(n1656), .B2(n1818), .ZN(n3534) );
  OAI22_X1 U949 ( .A1(n82), .A2(n1594), .B1(n1656), .B2(n1819), .ZN(n3533) );
  OAI22_X1 U950 ( .A1(n83), .A2(n1594), .B1(n1656), .B2(n1820), .ZN(n3532) );
  OAI22_X1 U951 ( .A1(n84), .A2(n1594), .B1(n1656), .B2(n1821), .ZN(n3531) );
  OAI22_X1 U952 ( .A1(n85), .A2(n1594), .B1(n1656), .B2(n1822), .ZN(n3530) );
  OAI22_X1 U953 ( .A1(n86), .A2(n1594), .B1(n1656), .B2(n1823), .ZN(n3529) );
  OAI22_X1 U954 ( .A1(n87), .A2(n1594), .B1(n1656), .B2(n1824), .ZN(n3528) );
  OAI22_X1 U955 ( .A1(n88), .A2(n1594), .B1(n1656), .B2(n1825), .ZN(n3527) );
  OAI22_X1 U956 ( .A1(n89), .A2(n1699), .B1(n1698), .B2(n1826), .ZN(n3526) );
  OAI22_X1 U957 ( .A1(n90), .A2(n1699), .B1(n1656), .B2(n1827), .ZN(n3525) );
  OAI22_X1 U958 ( .A1(n91), .A2(n1699), .B1(n1656), .B2(n1828), .ZN(n3524) );
  OAI22_X1 U959 ( .A1(n92), .A2(n1699), .B1(n1656), .B2(n1829), .ZN(n3523) );
  OAI22_X1 U960 ( .A1(n93), .A2(n1699), .B1(n1698), .B2(n1830), .ZN(n3522) );
  OAI22_X1 U961 ( .A1(n94), .A2(n1699), .B1(n1698), .B2(n1831), .ZN(n3521) );
  OAI22_X1 U962 ( .A1(n95), .A2(n1594), .B1(n1656), .B2(n1832), .ZN(n3520) );
  OAI22_X1 U963 ( .A1(n96), .A2(n1594), .B1(n1656), .B2(n1833), .ZN(n3519) );
  NAND2_X1 U964 ( .A1(n1714), .A2(n1788), .ZN(n1700) );
  OAI22_X1 U965 ( .A1(n97), .A2(n1593), .B1(n1701), .B2(n1802), .ZN(n3518) );
  OAI22_X1 U966 ( .A1(n98), .A2(n1593), .B1(n1701), .B2(n1803), .ZN(n3517) );
  OAI22_X1 U967 ( .A1(n99), .A2(n1593), .B1(n1701), .B2(n1804), .ZN(n3516) );
  OAI22_X1 U968 ( .A1(n100), .A2(n1593), .B1(n1701), .B2(n1805), .ZN(n3515) );
  OAI22_X1 U969 ( .A1(n101), .A2(n1593), .B1(n1701), .B2(n1806), .ZN(n3514) );
  OAI22_X1 U970 ( .A1(n102), .A2(n1593), .B1(n1701), .B2(n1807), .ZN(n3513) );
  OAI22_X1 U971 ( .A1(n103), .A2(n1593), .B1(n1701), .B2(n1808), .ZN(n3512) );
  OAI22_X1 U972 ( .A1(n104), .A2(n1593), .B1(n1701), .B2(n1809), .ZN(n3511) );
  OAI22_X1 U973 ( .A1(n105), .A2(n1593), .B1(n1701), .B2(n1810), .ZN(n3510) );
  OAI22_X1 U974 ( .A1(n106), .A2(n1593), .B1(n1701), .B2(n1811), .ZN(n3509) );
  OAI22_X1 U975 ( .A1(n107), .A2(n1593), .B1(n1701), .B2(n1812), .ZN(n3508) );
  OAI22_X1 U976 ( .A1(n108), .A2(n1593), .B1(n1701), .B2(n1813), .ZN(n3507) );
  OAI22_X1 U977 ( .A1(n109), .A2(n1593), .B1(n1657), .B2(n1814), .ZN(n3506) );
  OAI22_X1 U978 ( .A1(n110), .A2(n1593), .B1(n1657), .B2(n1815), .ZN(n3505) );
  OAI22_X1 U979 ( .A1(n111), .A2(n1593), .B1(n1657), .B2(n1816), .ZN(n3504) );
  OAI22_X1 U980 ( .A1(n112), .A2(n1593), .B1(n1657), .B2(n1817), .ZN(n3503) );
  OAI22_X1 U981 ( .A1(n113), .A2(n1593), .B1(n1657), .B2(n1818), .ZN(n3502) );
  OAI22_X1 U982 ( .A1(n114), .A2(n1593), .B1(n1657), .B2(n1819), .ZN(n3501) );
  OAI22_X1 U983 ( .A1(n115), .A2(n1593), .B1(n1657), .B2(n1820), .ZN(n3500) );
  OAI22_X1 U984 ( .A1(n116), .A2(n1593), .B1(n1657), .B2(n1821), .ZN(n3499) );
  OAI22_X1 U985 ( .A1(n117), .A2(n1593), .B1(n1657), .B2(n1822), .ZN(n3498) );
  OAI22_X1 U986 ( .A1(n118), .A2(n1593), .B1(n1657), .B2(n1823), .ZN(n3497) );
  OAI22_X1 U987 ( .A1(n119), .A2(n1593), .B1(n1657), .B2(n1824), .ZN(n3496) );
  OAI22_X1 U988 ( .A1(n120), .A2(n1593), .B1(n1657), .B2(n1825), .ZN(n3495) );
  OAI22_X1 U989 ( .A1(n121), .A2(n1702), .B1(n1701), .B2(n1826), .ZN(n3494) );
  OAI22_X1 U990 ( .A1(n122), .A2(n1702), .B1(n1657), .B2(n1827), .ZN(n3493) );
  OAI22_X1 U991 ( .A1(n123), .A2(n1702), .B1(n1657), .B2(n1828), .ZN(n3492) );
  OAI22_X1 U992 ( .A1(n124), .A2(n1702), .B1(n1657), .B2(n1829), .ZN(n3491) );
  OAI22_X1 U993 ( .A1(n125), .A2(n1702), .B1(n1701), .B2(n1830), .ZN(n3490) );
  OAI22_X1 U994 ( .A1(n126), .A2(n1702), .B1(n1701), .B2(n1831), .ZN(n3489) );
  OAI22_X1 U995 ( .A1(n127), .A2(n1593), .B1(n1657), .B2(n1832), .ZN(n3488) );
  OAI22_X1 U996 ( .A1(n128), .A2(n1593), .B1(n1657), .B2(n1833), .ZN(n3487) );
  NAND2_X1 U997 ( .A1(n1714), .A2(n1792), .ZN(n1704) );
  OAI22_X1 U998 ( .A1(n129), .A2(n1599), .B1(n1705), .B2(n1802), .ZN(n3486) );
  OAI22_X1 U999 ( .A1(n130), .A2(n1599), .B1(n1705), .B2(n1803), .ZN(n3485) );
  OAI22_X1 U1000 ( .A1(n131), .A2(n1599), .B1(n1705), .B2(n1804), .ZN(n3484)
         );
  OAI22_X1 U1001 ( .A1(n132), .A2(n1599), .B1(n1705), .B2(n1805), .ZN(n3483)
         );
  OAI22_X1 U1002 ( .A1(n133), .A2(n1599), .B1(n1705), .B2(n1806), .ZN(n3482)
         );
  OAI22_X1 U1003 ( .A1(n134), .A2(n1599), .B1(n1705), .B2(n1807), .ZN(n3481)
         );
  OAI22_X1 U1004 ( .A1(n135), .A2(n1599), .B1(n1705), .B2(n1808), .ZN(n3480)
         );
  OAI22_X1 U1005 ( .A1(n136), .A2(n1599), .B1(n1705), .B2(n1809), .ZN(n3479)
         );
  OAI22_X1 U1006 ( .A1(n137), .A2(n1599), .B1(n1705), .B2(n1810), .ZN(n3478)
         );
  OAI22_X1 U1007 ( .A1(n138), .A2(n1599), .B1(n1705), .B2(n1811), .ZN(n3477)
         );
  OAI22_X1 U1008 ( .A1(n139), .A2(n1599), .B1(n1705), .B2(n1812), .ZN(n3476)
         );
  OAI22_X1 U1009 ( .A1(n140), .A2(n1599), .B1(n1705), .B2(n1813), .ZN(n3475)
         );
  OAI22_X1 U1010 ( .A1(n141), .A2(n1599), .B1(n1658), .B2(n1814), .ZN(n3474)
         );
  OAI22_X1 U1011 ( .A1(n142), .A2(n1599), .B1(n1658), .B2(n1815), .ZN(n3473)
         );
  OAI22_X1 U1012 ( .A1(n143), .A2(n1599), .B1(n1658), .B2(n1816), .ZN(n3472)
         );
  OAI22_X1 U1013 ( .A1(n144), .A2(n1599), .B1(n1658), .B2(n1817), .ZN(n3471)
         );
  OAI22_X1 U1014 ( .A1(n145), .A2(n1599), .B1(n1658), .B2(n1818), .ZN(n3470)
         );
  OAI22_X1 U1015 ( .A1(n146), .A2(n1599), .B1(n1658), .B2(n1819), .ZN(n3469)
         );
  OAI22_X1 U1016 ( .A1(n147), .A2(n1599), .B1(n1658), .B2(n1820), .ZN(n3468)
         );
  OAI22_X1 U1017 ( .A1(n148), .A2(n1599), .B1(n1658), .B2(n1821), .ZN(n3467)
         );
  OAI22_X1 U1018 ( .A1(n149), .A2(n1599), .B1(n1658), .B2(n1822), .ZN(n3466)
         );
  OAI22_X1 U1019 ( .A1(n150), .A2(n1599), .B1(n1658), .B2(n1823), .ZN(n3465)
         );
  OAI22_X1 U1020 ( .A1(n151), .A2(n1599), .B1(n1658), .B2(n1824), .ZN(n3464)
         );
  OAI22_X1 U1021 ( .A1(n152), .A2(n1599), .B1(n1658), .B2(n1825), .ZN(n3463)
         );
  OAI22_X1 U1022 ( .A1(n153), .A2(n1706), .B1(n1705), .B2(n1826), .ZN(n3462)
         );
  OAI22_X1 U1023 ( .A1(n154), .A2(n1706), .B1(n1658), .B2(n1827), .ZN(n3461)
         );
  OAI22_X1 U1024 ( .A1(n155), .A2(n1706), .B1(n1658), .B2(n1828), .ZN(n3460)
         );
  OAI22_X1 U1025 ( .A1(n156), .A2(n1706), .B1(n1658), .B2(n1829), .ZN(n3459)
         );
  OAI22_X1 U1026 ( .A1(n157), .A2(n1706), .B1(n1705), .B2(n1830), .ZN(n3458)
         );
  OAI22_X1 U1027 ( .A1(n158), .A2(n1706), .B1(n1705), .B2(n1831), .ZN(n3457)
         );
  OAI22_X1 U1028 ( .A1(n159), .A2(n1599), .B1(n1658), .B2(n1832), .ZN(n3456)
         );
  OAI22_X1 U1029 ( .A1(n160), .A2(n1599), .B1(n1658), .B2(n1833), .ZN(n3455)
         );
  NAND2_X1 U1030 ( .A1(n1714), .A2(n1796), .ZN(n1708) );
  OAI22_X1 U1031 ( .A1(n161), .A2(n1588), .B1(n1709), .B2(n1802), .ZN(n3454)
         );
  OAI22_X1 U1032 ( .A1(n162), .A2(n1588), .B1(n1709), .B2(n1803), .ZN(n3453)
         );
  OAI22_X1 U1033 ( .A1(n163), .A2(n1588), .B1(n1709), .B2(n1804), .ZN(n3452)
         );
  OAI22_X1 U1034 ( .A1(n164), .A2(n1588), .B1(n1709), .B2(n1805), .ZN(n3451)
         );
  OAI22_X1 U1035 ( .A1(n165), .A2(n1588), .B1(n1709), .B2(n1806), .ZN(n3450)
         );
  OAI22_X1 U1036 ( .A1(n166), .A2(n1588), .B1(n1709), .B2(n1807), .ZN(n3449)
         );
  OAI22_X1 U1037 ( .A1(n167), .A2(n1588), .B1(n1709), .B2(n1808), .ZN(n3448)
         );
  OAI22_X1 U1038 ( .A1(n168), .A2(n1588), .B1(n1709), .B2(n1809), .ZN(n3447)
         );
  OAI22_X1 U1039 ( .A1(n169), .A2(n1588), .B1(n1709), .B2(n1810), .ZN(n3446)
         );
  OAI22_X1 U1040 ( .A1(n170), .A2(n1588), .B1(n1709), .B2(n1811), .ZN(n3445)
         );
  OAI22_X1 U1041 ( .A1(n171), .A2(n1588), .B1(n1709), .B2(n1812), .ZN(n3444)
         );
  OAI22_X1 U1042 ( .A1(n172), .A2(n1588), .B1(n1709), .B2(n1813), .ZN(n3443)
         );
  OAI22_X1 U1043 ( .A1(n173), .A2(n1588), .B1(n1659), .B2(n1814), .ZN(n3442)
         );
  OAI22_X1 U1044 ( .A1(n174), .A2(n1588), .B1(n1659), .B2(n1815), .ZN(n3441)
         );
  OAI22_X1 U1045 ( .A1(n175), .A2(n1588), .B1(n1659), .B2(n1816), .ZN(n3440)
         );
  OAI22_X1 U1046 ( .A1(n176), .A2(n1588), .B1(n1659), .B2(n1817), .ZN(n3439)
         );
  OAI22_X1 U1047 ( .A1(n177), .A2(n1588), .B1(n1659), .B2(n1818), .ZN(n3438)
         );
  OAI22_X1 U1048 ( .A1(n178), .A2(n1588), .B1(n1659), .B2(n1819), .ZN(n3437)
         );
  OAI22_X1 U1049 ( .A1(n179), .A2(n1588), .B1(n1659), .B2(n1820), .ZN(n3436)
         );
  OAI22_X1 U1050 ( .A1(n180), .A2(n1588), .B1(n1659), .B2(n1821), .ZN(n3435)
         );
  OAI22_X1 U1051 ( .A1(n181), .A2(n1588), .B1(n1659), .B2(n1822), .ZN(n3434)
         );
  OAI22_X1 U1052 ( .A1(n182), .A2(n1588), .B1(n1659), .B2(n1823), .ZN(n3433)
         );
  OAI22_X1 U1053 ( .A1(n183), .A2(n1588), .B1(n1659), .B2(n1824), .ZN(n3432)
         );
  OAI22_X1 U1054 ( .A1(n184), .A2(n1588), .B1(n1659), .B2(n1825), .ZN(n3431)
         );
  OAI22_X1 U1055 ( .A1(n185), .A2(n1710), .B1(n1709), .B2(n1826), .ZN(n3430)
         );
  OAI22_X1 U1056 ( .A1(n186), .A2(n1710), .B1(n1659), .B2(n1827), .ZN(n3429)
         );
  OAI22_X1 U1057 ( .A1(n187), .A2(n1710), .B1(n1659), .B2(n1828), .ZN(n3428)
         );
  OAI22_X1 U1058 ( .A1(n188), .A2(n1710), .B1(n1659), .B2(n1829), .ZN(n3427)
         );
  OAI22_X1 U1059 ( .A1(n189), .A2(n1710), .B1(n1709), .B2(n1830), .ZN(n3426)
         );
  OAI22_X1 U1060 ( .A1(n190), .A2(n1710), .B1(n1709), .B2(n1831), .ZN(n3425)
         );
  OAI22_X1 U1061 ( .A1(n191), .A2(n1588), .B1(n1659), .B2(n1832), .ZN(n3424)
         );
  OAI22_X1 U1062 ( .A1(n192), .A2(n1588), .B1(n1659), .B2(n1833), .ZN(n3423)
         );
  NAND2_X1 U1063 ( .A1(n1714), .A2(n1801), .ZN(n1713) );
  OAI22_X1 U1064 ( .A1(n193), .A2(n1595), .B1(n1715), .B2(n1802), .ZN(n3422)
         );
  OAI22_X1 U1065 ( .A1(n194), .A2(n1595), .B1(n1715), .B2(n1803), .ZN(n3421)
         );
  OAI22_X1 U1066 ( .A1(n195), .A2(n1595), .B1(n1715), .B2(n1804), .ZN(n3420)
         );
  OAI22_X1 U1067 ( .A1(n196), .A2(n1595), .B1(n1715), .B2(n1805), .ZN(n3419)
         );
  OAI22_X1 U1068 ( .A1(n197), .A2(n1595), .B1(n1715), .B2(n1806), .ZN(n3418)
         );
  OAI22_X1 U1069 ( .A1(n198), .A2(n1595), .B1(n1715), .B2(n1807), .ZN(n3417)
         );
  OAI22_X1 U1070 ( .A1(n199), .A2(n1595), .B1(n1715), .B2(n1808), .ZN(n3416)
         );
  OAI22_X1 U1071 ( .A1(n200), .A2(n1595), .B1(n1715), .B2(n1809), .ZN(n3415)
         );
  OAI22_X1 U1072 ( .A1(n201), .A2(n1595), .B1(n1715), .B2(n1810), .ZN(n3414)
         );
  OAI22_X1 U1073 ( .A1(n202), .A2(n1595), .B1(n1715), .B2(n1811), .ZN(n3413)
         );
  OAI22_X1 U1074 ( .A1(n203), .A2(n1595), .B1(n1715), .B2(n1812), .ZN(n3412)
         );
  OAI22_X1 U1075 ( .A1(n204), .A2(n1595), .B1(n1715), .B2(n1813), .ZN(n3411)
         );
  OAI22_X1 U1076 ( .A1(n205), .A2(n1595), .B1(n1660), .B2(n1814), .ZN(n3410)
         );
  OAI22_X1 U1077 ( .A1(n206), .A2(n1595), .B1(n1660), .B2(n1815), .ZN(n3409)
         );
  OAI22_X1 U1078 ( .A1(n207), .A2(n1595), .B1(n1660), .B2(n1816), .ZN(n3408)
         );
  OAI22_X1 U1079 ( .A1(n208), .A2(n1595), .B1(n1660), .B2(n1817), .ZN(n3407)
         );
  OAI22_X1 U1080 ( .A1(n209), .A2(n1595), .B1(n1660), .B2(n1818), .ZN(n3406)
         );
  OAI22_X1 U1081 ( .A1(n210), .A2(n1595), .B1(n1660), .B2(n1819), .ZN(n3405)
         );
  OAI22_X1 U1082 ( .A1(n211), .A2(n1595), .B1(n1660), .B2(n1820), .ZN(n3404)
         );
  OAI22_X1 U1083 ( .A1(n212), .A2(n1595), .B1(n1660), .B2(n1821), .ZN(n3403)
         );
  OAI22_X1 U1084 ( .A1(n213), .A2(n1595), .B1(n1660), .B2(n1822), .ZN(n3402)
         );
  OAI22_X1 U1085 ( .A1(n214), .A2(n1595), .B1(n1660), .B2(n1823), .ZN(n3401)
         );
  OAI22_X1 U1086 ( .A1(n215), .A2(n1595), .B1(n1660), .B2(n1824), .ZN(n3400)
         );
  OAI22_X1 U1087 ( .A1(n216), .A2(n1595), .B1(n1660), .B2(n1825), .ZN(n3399)
         );
  OAI22_X1 U1088 ( .A1(n217), .A2(n1716), .B1(n1715), .B2(n1826), .ZN(n3398)
         );
  OAI22_X1 U1089 ( .A1(n218), .A2(n1716), .B1(n1660), .B2(n1827), .ZN(n3397)
         );
  OAI22_X1 U1090 ( .A1(n219), .A2(n1716), .B1(n1660), .B2(n1828), .ZN(n3396)
         );
  OAI22_X1 U1091 ( .A1(n220), .A2(n1716), .B1(n1660), .B2(n1829), .ZN(n3395)
         );
  OAI22_X1 U1092 ( .A1(n221), .A2(n1716), .B1(n1715), .B2(n1830), .ZN(n3394)
         );
  OAI22_X1 U1093 ( .A1(n222), .A2(n1716), .B1(n1715), .B2(n1831), .ZN(n3393)
         );
  OAI22_X1 U1094 ( .A1(n223), .A2(n1595), .B1(n1660), .B2(n1832), .ZN(n3392)
         );
  OAI22_X1 U1095 ( .A1(n224), .A2(n1595), .B1(n1660), .B2(n1833), .ZN(n3391)
         );
  NAND2_X1 U1096 ( .A1(n1772), .A2(n1740), .ZN(n1717) );
  OAI22_X1 U1097 ( .A1(n225), .A2(n1614), .B1(n1719), .B2(n1802), .ZN(n3390)
         );
  OAI22_X1 U1098 ( .A1(n226), .A2(n1614), .B1(n1719), .B2(n1803), .ZN(n3389)
         );
  OAI22_X1 U1099 ( .A1(n227), .A2(n1614), .B1(n1719), .B2(n1804), .ZN(n3388)
         );
  OAI22_X1 U1100 ( .A1(n228), .A2(n1614), .B1(n1719), .B2(n1805), .ZN(n3387)
         );
  OAI22_X1 U1101 ( .A1(n229), .A2(n1614), .B1(n1719), .B2(n1806), .ZN(n3386)
         );
  OAI22_X1 U1102 ( .A1(n230), .A2(n1614), .B1(n1719), .B2(n1807), .ZN(n3385)
         );
  OAI22_X1 U1103 ( .A1(n231), .A2(n1614), .B1(n1719), .B2(n1808), .ZN(n3384)
         );
  OAI22_X1 U1104 ( .A1(n232), .A2(n1614), .B1(n1719), .B2(n1809), .ZN(n3383)
         );
  OAI22_X1 U1105 ( .A1(n233), .A2(n1614), .B1(n1719), .B2(n1810), .ZN(n3382)
         );
  OAI22_X1 U1106 ( .A1(n234), .A2(n1614), .B1(n1719), .B2(n1811), .ZN(n3381)
         );
  OAI22_X1 U1107 ( .A1(n235), .A2(n1614), .B1(n1719), .B2(n1812), .ZN(n3380)
         );
  OAI22_X1 U1108 ( .A1(n236), .A2(n1614), .B1(n1719), .B2(n1813), .ZN(n3379)
         );
  OAI22_X1 U1109 ( .A1(n237), .A2(n1614), .B1(n1719), .B2(n1814), .ZN(n3378)
         );
  OAI22_X1 U1110 ( .A1(n238), .A2(n1614), .B1(n1719), .B2(n1815), .ZN(n3377)
         );
  OAI22_X1 U1111 ( .A1(n239), .A2(n1614), .B1(n1719), .B2(n1816), .ZN(n3376)
         );
  OAI22_X1 U1112 ( .A1(n240), .A2(n1614), .B1(n1719), .B2(n1817), .ZN(n3375)
         );
  OAI22_X1 U1113 ( .A1(n241), .A2(n1614), .B1(n1719), .B2(n1818), .ZN(n3374)
         );
  OAI22_X1 U1114 ( .A1(n242), .A2(n1614), .B1(n1719), .B2(n1819), .ZN(n3373)
         );
  OAI22_X1 U1115 ( .A1(n243), .A2(n1614), .B1(n1719), .B2(n1820), .ZN(n3372)
         );
  OAI22_X1 U1116 ( .A1(n244), .A2(n1614), .B1(n1719), .B2(n1821), .ZN(n3371)
         );
  OAI22_X1 U1117 ( .A1(n245), .A2(n1614), .B1(n1719), .B2(n1822), .ZN(n3370)
         );
  OAI22_X1 U1118 ( .A1(n246), .A2(n1614), .B1(n1719), .B2(n1823), .ZN(n3369)
         );
  OAI22_X1 U1119 ( .A1(n247), .A2(n1614), .B1(n1719), .B2(n1824), .ZN(n3368)
         );
  OAI22_X1 U1120 ( .A1(n248), .A2(n1614), .B1(n1719), .B2(n1825), .ZN(n3367)
         );
  OAI22_X1 U1121 ( .A1(n249), .A2(n1720), .B1(n1719), .B2(n1826), .ZN(n3366)
         );
  OAI22_X1 U1122 ( .A1(n250), .A2(n1720), .B1(n1719), .B2(n1827), .ZN(n3365)
         );
  OAI22_X1 U1123 ( .A1(n251), .A2(n1720), .B1(n1719), .B2(n1828), .ZN(n3364)
         );
  OAI22_X1 U1124 ( .A1(n252), .A2(n1720), .B1(n1719), .B2(n1829), .ZN(n3363)
         );
  OAI22_X1 U1125 ( .A1(n253), .A2(n1720), .B1(n1719), .B2(n1830), .ZN(n3362)
         );
  OAI22_X1 U1126 ( .A1(n254), .A2(n1720), .B1(n1719), .B2(n1831), .ZN(n3361)
         );
  OAI22_X1 U1127 ( .A1(n255), .A2(n1614), .B1(n1719), .B2(n1832), .ZN(n3360)
         );
  OAI22_X1 U1128 ( .A1(n256), .A2(n1614), .B1(n1719), .B2(n1833), .ZN(n3359)
         );
  NAND2_X1 U1129 ( .A1(n1776), .A2(n1740), .ZN(n1721) );
  OAI22_X1 U1130 ( .A1(n257), .A2(n1598), .B1(n1722), .B2(n1802), .ZN(n3358)
         );
  OAI22_X1 U1131 ( .A1(n258), .A2(n1598), .B1(n1722), .B2(n1803), .ZN(n3357)
         );
  OAI22_X1 U1132 ( .A1(n259), .A2(n1598), .B1(n1722), .B2(n1804), .ZN(n3356)
         );
  OAI22_X1 U1133 ( .A1(n260), .A2(n1598), .B1(n1722), .B2(n1805), .ZN(n3355)
         );
  OAI22_X1 U1134 ( .A1(n261), .A2(n1598), .B1(n1722), .B2(n1806), .ZN(n3354)
         );
  OAI22_X1 U1135 ( .A1(n262), .A2(n1598), .B1(n1722), .B2(n1807), .ZN(n3353)
         );
  OAI22_X1 U1136 ( .A1(n263), .A2(n1598), .B1(n1722), .B2(n1808), .ZN(n3352)
         );
  OAI22_X1 U1137 ( .A1(n264), .A2(n1598), .B1(n1722), .B2(n1809), .ZN(n3351)
         );
  OAI22_X1 U1138 ( .A1(n265), .A2(n1598), .B1(n1722), .B2(n1810), .ZN(n3350)
         );
  OAI22_X1 U1139 ( .A1(n266), .A2(n1598), .B1(n1722), .B2(n1811), .ZN(n3349)
         );
  OAI22_X1 U1140 ( .A1(n267), .A2(n1598), .B1(n1722), .B2(n1812), .ZN(n3348)
         );
  OAI22_X1 U1141 ( .A1(n268), .A2(n1598), .B1(n1722), .B2(n1813), .ZN(n3347)
         );
  OAI22_X1 U1142 ( .A1(n269), .A2(n1598), .B1(n1661), .B2(n1814), .ZN(n3346)
         );
  OAI22_X1 U1143 ( .A1(n270), .A2(n1598), .B1(n1661), .B2(n1815), .ZN(n3345)
         );
  OAI22_X1 U1144 ( .A1(n271), .A2(n1598), .B1(n1661), .B2(n1816), .ZN(n3344)
         );
  OAI22_X1 U1145 ( .A1(n272), .A2(n1598), .B1(n1661), .B2(n1817), .ZN(n3343)
         );
  OAI22_X1 U1146 ( .A1(n273), .A2(n1598), .B1(n1661), .B2(n1818), .ZN(n3342)
         );
  OAI22_X1 U1147 ( .A1(n274), .A2(n1598), .B1(n1661), .B2(n1819), .ZN(n3341)
         );
  OAI22_X1 U1148 ( .A1(n275), .A2(n1598), .B1(n1661), .B2(n1820), .ZN(n3340)
         );
  OAI22_X1 U1149 ( .A1(n276), .A2(n1598), .B1(n1661), .B2(n1821), .ZN(n3339)
         );
  OAI22_X1 U1150 ( .A1(n277), .A2(n1598), .B1(n1661), .B2(n1822), .ZN(n3338)
         );
  OAI22_X1 U1151 ( .A1(n278), .A2(n1598), .B1(n1661), .B2(n1823), .ZN(n3337)
         );
  OAI22_X1 U1152 ( .A1(n279), .A2(n1598), .B1(n1661), .B2(n1824), .ZN(n3336)
         );
  OAI22_X1 U1153 ( .A1(n280), .A2(n1598), .B1(n1661), .B2(n1825), .ZN(n3335)
         );
  OAI22_X1 U1154 ( .A1(n281), .A2(n1723), .B1(n1661), .B2(n1826), .ZN(n3334)
         );
  OAI22_X1 U1155 ( .A1(n282), .A2(n1723), .B1(n1661), .B2(n1827), .ZN(n3333)
         );
  OAI22_X1 U1156 ( .A1(n283), .A2(n1723), .B1(n1661), .B2(n1828), .ZN(n3332)
         );
  OAI22_X1 U1157 ( .A1(n284), .A2(n1723), .B1(n1661), .B2(n1829), .ZN(n3331)
         );
  OAI22_X1 U1158 ( .A1(n285), .A2(n1723), .B1(n1722), .B2(n1830), .ZN(n3330)
         );
  OAI22_X1 U1159 ( .A1(n286), .A2(n1723), .B1(n1722), .B2(n1831), .ZN(n3329)
         );
  OAI22_X1 U1160 ( .A1(n287), .A2(n1598), .B1(n1722), .B2(n1832), .ZN(n3328)
         );
  OAI22_X1 U1161 ( .A1(n288), .A2(n1598), .B1(n1722), .B2(n1833), .ZN(n3327)
         );
  NAND2_X1 U1162 ( .A1(n1780), .A2(n1740), .ZN(n1724) );
  OAI22_X1 U1163 ( .A1(n289), .A2(n1590), .B1(n1725), .B2(n1802), .ZN(n3326)
         );
  OAI22_X1 U1164 ( .A1(n290), .A2(n1590), .B1(n1725), .B2(n1803), .ZN(n3325)
         );
  OAI22_X1 U1165 ( .A1(n291), .A2(n1590), .B1(n1725), .B2(n1804), .ZN(n3324)
         );
  OAI22_X1 U1166 ( .A1(n292), .A2(n1590), .B1(n1725), .B2(n1805), .ZN(n3323)
         );
  OAI22_X1 U1167 ( .A1(n293), .A2(n1590), .B1(n1725), .B2(n1806), .ZN(n3322)
         );
  OAI22_X1 U1168 ( .A1(n294), .A2(n1590), .B1(n1725), .B2(n1807), .ZN(n3321)
         );
  OAI22_X1 U1169 ( .A1(n295), .A2(n1590), .B1(n1725), .B2(n1808), .ZN(n3320)
         );
  OAI22_X1 U1170 ( .A1(n296), .A2(n1590), .B1(n1725), .B2(n1809), .ZN(n3319)
         );
  OAI22_X1 U1171 ( .A1(n297), .A2(n1590), .B1(n1725), .B2(n1810), .ZN(n3318)
         );
  OAI22_X1 U1172 ( .A1(n298), .A2(n1590), .B1(n1725), .B2(n1811), .ZN(n3317)
         );
  OAI22_X1 U1173 ( .A1(n299), .A2(n1590), .B1(n1725), .B2(n1812), .ZN(n3316)
         );
  OAI22_X1 U1174 ( .A1(n300), .A2(n1590), .B1(n1725), .B2(n1813), .ZN(n3315)
         );
  OAI22_X1 U1175 ( .A1(n301), .A2(n1590), .B1(n1662), .B2(n1814), .ZN(n3314)
         );
  OAI22_X1 U1176 ( .A1(n302), .A2(n1590), .B1(n1662), .B2(n1815), .ZN(n3313)
         );
  OAI22_X1 U1177 ( .A1(n303), .A2(n1590), .B1(n1662), .B2(n1816), .ZN(n3312)
         );
  OAI22_X1 U1178 ( .A1(n304), .A2(n1590), .B1(n1662), .B2(n1817), .ZN(n3311)
         );
  OAI22_X1 U1179 ( .A1(n305), .A2(n1590), .B1(n1662), .B2(n1818), .ZN(n3310)
         );
  OAI22_X1 U1180 ( .A1(n306), .A2(n1590), .B1(n1662), .B2(n1819), .ZN(n3309)
         );
  OAI22_X1 U1181 ( .A1(n307), .A2(n1590), .B1(n1662), .B2(n1820), .ZN(n3308)
         );
  OAI22_X1 U1182 ( .A1(n308), .A2(n1590), .B1(n1662), .B2(n1821), .ZN(n3307)
         );
  OAI22_X1 U1183 ( .A1(n309), .A2(n1590), .B1(n1662), .B2(n1822), .ZN(n3306)
         );
  OAI22_X1 U1184 ( .A1(n310), .A2(n1590), .B1(n1662), .B2(n1823), .ZN(n3305)
         );
  OAI22_X1 U1185 ( .A1(n311), .A2(n1590), .B1(n1662), .B2(n1824), .ZN(n3304)
         );
  OAI22_X1 U1186 ( .A1(n312), .A2(n1590), .B1(n1662), .B2(n1825), .ZN(n3303)
         );
  OAI22_X1 U1187 ( .A1(n313), .A2(n1726), .B1(n1662), .B2(n1826), .ZN(n3302)
         );
  OAI22_X1 U1188 ( .A1(n314), .A2(n1726), .B1(n1662), .B2(n1827), .ZN(n3301)
         );
  OAI22_X1 U1189 ( .A1(n315), .A2(n1726), .B1(n1662), .B2(n1828), .ZN(n3300)
         );
  OAI22_X1 U1190 ( .A1(n316), .A2(n1726), .B1(n1662), .B2(n1829), .ZN(n3299)
         );
  OAI22_X1 U1191 ( .A1(n317), .A2(n1726), .B1(n1725), .B2(n1830), .ZN(n3298)
         );
  OAI22_X1 U1192 ( .A1(n318), .A2(n1726), .B1(n1725), .B2(n1831), .ZN(n3297)
         );
  OAI22_X1 U1193 ( .A1(n319), .A2(n1590), .B1(n1725), .B2(n1832), .ZN(n3296)
         );
  OAI22_X1 U1194 ( .A1(n320), .A2(n1590), .B1(n1725), .B2(n1833), .ZN(n3295)
         );
  NAND2_X1 U1195 ( .A1(n1784), .A2(n1740), .ZN(n1727) );
  OAI22_X1 U1196 ( .A1(n321), .A2(n1597), .B1(n1728), .B2(n1802), .ZN(n3294)
         );
  OAI22_X1 U1197 ( .A1(n322), .A2(n1597), .B1(n1728), .B2(n1803), .ZN(n3293)
         );
  OAI22_X1 U1198 ( .A1(n323), .A2(n1597), .B1(n1728), .B2(n1804), .ZN(n3292)
         );
  OAI22_X1 U1199 ( .A1(n324), .A2(n1597), .B1(n1728), .B2(n1805), .ZN(n3291)
         );
  OAI22_X1 U1200 ( .A1(n325), .A2(n1597), .B1(n1728), .B2(n1806), .ZN(n3290)
         );
  OAI22_X1 U1201 ( .A1(n326), .A2(n1597), .B1(n1728), .B2(n1807), .ZN(n3289)
         );
  OAI22_X1 U1202 ( .A1(n327), .A2(n1597), .B1(n1728), .B2(n1808), .ZN(n3288)
         );
  OAI22_X1 U1203 ( .A1(n328), .A2(n1597), .B1(n1728), .B2(n1809), .ZN(n3287)
         );
  OAI22_X1 U1204 ( .A1(n329), .A2(n1597), .B1(n1728), .B2(n1810), .ZN(n3286)
         );
  OAI22_X1 U1205 ( .A1(n330), .A2(n1597), .B1(n1728), .B2(n1811), .ZN(n3285)
         );
  OAI22_X1 U1206 ( .A1(n331), .A2(n1597), .B1(n1728), .B2(n1812), .ZN(n3284)
         );
  OAI22_X1 U1207 ( .A1(n332), .A2(n1597), .B1(n1728), .B2(n1813), .ZN(n3283)
         );
  OAI22_X1 U1208 ( .A1(n333), .A2(n1597), .B1(n1663), .B2(n1814), .ZN(n3282)
         );
  OAI22_X1 U1209 ( .A1(n334), .A2(n1597), .B1(n1663), .B2(n1815), .ZN(n3281)
         );
  OAI22_X1 U1210 ( .A1(n335), .A2(n1597), .B1(n1663), .B2(n1816), .ZN(n3280)
         );
  OAI22_X1 U1211 ( .A1(n336), .A2(n1597), .B1(n1663), .B2(n1817), .ZN(n3279)
         );
  OAI22_X1 U1212 ( .A1(n337), .A2(n1597), .B1(n1663), .B2(n1818), .ZN(n3278)
         );
  OAI22_X1 U1213 ( .A1(n338), .A2(n1597), .B1(n1663), .B2(n1819), .ZN(n3277)
         );
  OAI22_X1 U1214 ( .A1(n339), .A2(n1597), .B1(n1663), .B2(n1820), .ZN(n3276)
         );
  OAI22_X1 U1215 ( .A1(n340), .A2(n1597), .B1(n1663), .B2(n1821), .ZN(n3275)
         );
  OAI22_X1 U1216 ( .A1(n341), .A2(n1597), .B1(n1663), .B2(n1822), .ZN(n3274)
         );
  OAI22_X1 U1217 ( .A1(n342), .A2(n1597), .B1(n1663), .B2(n1823), .ZN(n3273)
         );
  OAI22_X1 U1218 ( .A1(n343), .A2(n1597), .B1(n1663), .B2(n1824), .ZN(n3272)
         );
  OAI22_X1 U1219 ( .A1(n344), .A2(n1597), .B1(n1663), .B2(n1825), .ZN(n3271)
         );
  OAI22_X1 U1220 ( .A1(n345), .A2(n1729), .B1(n1663), .B2(n1826), .ZN(n3270)
         );
  OAI22_X1 U1221 ( .A1(n346), .A2(n1729), .B1(n1663), .B2(n1827), .ZN(n3269)
         );
  OAI22_X1 U1222 ( .A1(n347), .A2(n1729), .B1(n1663), .B2(n1828), .ZN(n3268)
         );
  OAI22_X1 U1223 ( .A1(n348), .A2(n1729), .B1(n1663), .B2(n1829), .ZN(n3267)
         );
  OAI22_X1 U1224 ( .A1(n349), .A2(n1729), .B1(n1728), .B2(n1830), .ZN(n3266)
         );
  OAI22_X1 U1225 ( .A1(n350), .A2(n1729), .B1(n1728), .B2(n1831), .ZN(n3265)
         );
  OAI22_X1 U1226 ( .A1(n351), .A2(n1597), .B1(n1728), .B2(n1832), .ZN(n3264)
         );
  OAI22_X1 U1227 ( .A1(n352), .A2(n1597), .B1(n1728), .B2(n1833), .ZN(n3263)
         );
  NAND2_X1 U1228 ( .A1(n1788), .A2(n1740), .ZN(n1730) );
  OAI22_X1 U1229 ( .A1(n353), .A2(n1611), .B1(n1731), .B2(n1802), .ZN(n3262)
         );
  OAI22_X1 U1230 ( .A1(n354), .A2(n1611), .B1(n1731), .B2(n1803), .ZN(n3261)
         );
  OAI22_X1 U1231 ( .A1(n355), .A2(n1611), .B1(n1731), .B2(n1804), .ZN(n3260)
         );
  OAI22_X1 U1232 ( .A1(n356), .A2(n1611), .B1(n1731), .B2(n1805), .ZN(n3259)
         );
  OAI22_X1 U1233 ( .A1(n357), .A2(n1611), .B1(n1731), .B2(n1806), .ZN(n3258)
         );
  OAI22_X1 U1234 ( .A1(n358), .A2(n1611), .B1(n1731), .B2(n1807), .ZN(n3257)
         );
  OAI22_X1 U1235 ( .A1(n359), .A2(n1611), .B1(n1731), .B2(n1808), .ZN(n3256)
         );
  OAI22_X1 U1236 ( .A1(n360), .A2(n1611), .B1(n1731), .B2(n1809), .ZN(n3255)
         );
  OAI22_X1 U1237 ( .A1(n361), .A2(n1611), .B1(n1731), .B2(n1810), .ZN(n3254)
         );
  OAI22_X1 U1238 ( .A1(n362), .A2(n1611), .B1(n1731), .B2(n1811), .ZN(n3253)
         );
  OAI22_X1 U1239 ( .A1(n363), .A2(n1611), .B1(n1731), .B2(n1812), .ZN(n3252)
         );
  OAI22_X1 U1240 ( .A1(n364), .A2(n1611), .B1(n1731), .B2(n1813), .ZN(n3251)
         );
  OAI22_X1 U1241 ( .A1(n365), .A2(n1611), .B1(n1664), .B2(n1814), .ZN(n3250)
         );
  OAI22_X1 U1242 ( .A1(n366), .A2(n1611), .B1(n1664), .B2(n1815), .ZN(n3249)
         );
  OAI22_X1 U1243 ( .A1(n367), .A2(n1611), .B1(n1664), .B2(n1816), .ZN(n3248)
         );
  OAI22_X1 U1244 ( .A1(n368), .A2(n1611), .B1(n1664), .B2(n1817), .ZN(n3247)
         );
  OAI22_X1 U1245 ( .A1(n369), .A2(n1611), .B1(n1664), .B2(n1818), .ZN(n3246)
         );
  OAI22_X1 U1246 ( .A1(n370), .A2(n1611), .B1(n1664), .B2(n1819), .ZN(n3245)
         );
  OAI22_X1 U1247 ( .A1(n371), .A2(n1611), .B1(n1664), .B2(n1820), .ZN(n3244)
         );
  OAI22_X1 U1248 ( .A1(n372), .A2(n1611), .B1(n1664), .B2(n1821), .ZN(n3243)
         );
  OAI22_X1 U1249 ( .A1(n373), .A2(n1611), .B1(n1664), .B2(n1822), .ZN(n3242)
         );
  OAI22_X1 U1250 ( .A1(n374), .A2(n1611), .B1(n1664), .B2(n1823), .ZN(n3241)
         );
  OAI22_X1 U1251 ( .A1(n375), .A2(n1611), .B1(n1664), .B2(n1824), .ZN(n3240)
         );
  OAI22_X1 U1252 ( .A1(n376), .A2(n1611), .B1(n1664), .B2(n1825), .ZN(n3239)
         );
  OAI22_X1 U1253 ( .A1(n377), .A2(n1732), .B1(n1664), .B2(n1826), .ZN(n3238)
         );
  OAI22_X1 U1254 ( .A1(n378), .A2(n1732), .B1(n1664), .B2(n1827), .ZN(n3237)
         );
  OAI22_X1 U1255 ( .A1(n379), .A2(n1732), .B1(n1664), .B2(n1828), .ZN(n3236)
         );
  OAI22_X1 U1256 ( .A1(n380), .A2(n1732), .B1(n1664), .B2(n1829), .ZN(n3235)
         );
  OAI22_X1 U1257 ( .A1(n381), .A2(n1732), .B1(n1731), .B2(n1830), .ZN(n3234)
         );
  OAI22_X1 U1258 ( .A1(n382), .A2(n1732), .B1(n1731), .B2(n1831), .ZN(n3233)
         );
  OAI22_X1 U1259 ( .A1(n383), .A2(n1611), .B1(n1731), .B2(n1832), .ZN(n3232)
         );
  OAI22_X1 U1260 ( .A1(n384), .A2(n1611), .B1(n1731), .B2(n1833), .ZN(n3231)
         );
  NAND2_X1 U1261 ( .A1(n1792), .A2(n1740), .ZN(n1733) );
  OAI22_X1 U1262 ( .A1(n385), .A2(n1604), .B1(n1734), .B2(n1802), .ZN(n3230)
         );
  OAI22_X1 U1263 ( .A1(n386), .A2(n1604), .B1(n1734), .B2(n1803), .ZN(n3229)
         );
  OAI22_X1 U1264 ( .A1(n387), .A2(n1604), .B1(n1734), .B2(n1804), .ZN(n3228)
         );
  OAI22_X1 U1265 ( .A1(n388), .A2(n1604), .B1(n1734), .B2(n1805), .ZN(n3227)
         );
  OAI22_X1 U1266 ( .A1(n389), .A2(n1604), .B1(n1734), .B2(n1806), .ZN(n3226)
         );
  OAI22_X1 U1267 ( .A1(n390), .A2(n1604), .B1(n1734), .B2(n1807), .ZN(n3225)
         );
  OAI22_X1 U1268 ( .A1(n391), .A2(n1604), .B1(n1734), .B2(n1808), .ZN(n3224)
         );
  OAI22_X1 U1269 ( .A1(n392), .A2(n1604), .B1(n1734), .B2(n1809), .ZN(n3223)
         );
  OAI22_X1 U1270 ( .A1(n393), .A2(n1604), .B1(n1734), .B2(n1810), .ZN(n3222)
         );
  OAI22_X1 U1271 ( .A1(n394), .A2(n1604), .B1(n1734), .B2(n1811), .ZN(n3221)
         );
  OAI22_X1 U1272 ( .A1(n395), .A2(n1604), .B1(n1734), .B2(n1812), .ZN(n3220)
         );
  OAI22_X1 U1273 ( .A1(n396), .A2(n1604), .B1(n1734), .B2(n1813), .ZN(n3219)
         );
  OAI22_X1 U1274 ( .A1(n397), .A2(n1604), .B1(n1665), .B2(n1814), .ZN(n3218)
         );
  OAI22_X1 U1275 ( .A1(n398), .A2(n1604), .B1(n1665), .B2(n1815), .ZN(n3217)
         );
  OAI22_X1 U1276 ( .A1(n399), .A2(n1604), .B1(n1665), .B2(n1816), .ZN(n3216)
         );
  OAI22_X1 U1277 ( .A1(n400), .A2(n1604), .B1(n1665), .B2(n1817), .ZN(n3215)
         );
  OAI22_X1 U1278 ( .A1(n401), .A2(n1604), .B1(n1665), .B2(n1818), .ZN(n3214)
         );
  OAI22_X1 U1279 ( .A1(n402), .A2(n1604), .B1(n1665), .B2(n1819), .ZN(n3213)
         );
  OAI22_X1 U1280 ( .A1(n403), .A2(n1604), .B1(n1665), .B2(n1820), .ZN(n3212)
         );
  OAI22_X1 U1281 ( .A1(n404), .A2(n1604), .B1(n1665), .B2(n1821), .ZN(n3211)
         );
  OAI22_X1 U1282 ( .A1(n405), .A2(n1604), .B1(n1665), .B2(n1822), .ZN(n3210)
         );
  OAI22_X1 U1283 ( .A1(n406), .A2(n1604), .B1(n1665), .B2(n1823), .ZN(n3209)
         );
  OAI22_X1 U1284 ( .A1(n407), .A2(n1604), .B1(n1665), .B2(n1824), .ZN(n3208)
         );
  OAI22_X1 U1285 ( .A1(n408), .A2(n1604), .B1(n1665), .B2(n1825), .ZN(n3207)
         );
  OAI22_X1 U1286 ( .A1(n409), .A2(n1735), .B1(n1665), .B2(n1826), .ZN(n3206)
         );
  OAI22_X1 U1287 ( .A1(n410), .A2(n1735), .B1(n1665), .B2(n1827), .ZN(n3205)
         );
  OAI22_X1 U1288 ( .A1(n411), .A2(n1604), .B1(n1665), .B2(n1828), .ZN(n3204)
         );
  OAI22_X1 U1289 ( .A1(n412), .A2(n1735), .B1(n1665), .B2(n1829), .ZN(n3203)
         );
  OAI22_X1 U1290 ( .A1(n413), .A2(n1735), .B1(n1734), .B2(n1830), .ZN(n3202)
         );
  OAI22_X1 U1291 ( .A1(n414), .A2(n1735), .B1(n1734), .B2(n1831), .ZN(n3201)
         );
  OAI22_X1 U1292 ( .A1(n415), .A2(n1735), .B1(n1734), .B2(n1832), .ZN(n3200)
         );
  OAI22_X1 U1293 ( .A1(n416), .A2(n1604), .B1(n1734), .B2(n1833), .ZN(n3199)
         );
  NAND2_X1 U1294 ( .A1(n1796), .A2(n1740), .ZN(n1736) );
  OAI22_X1 U1295 ( .A1(n417), .A2(n1583), .B1(n1737), .B2(n1802), .ZN(n3198)
         );
  OAI22_X1 U1296 ( .A1(n418), .A2(n1583), .B1(n1737), .B2(n1803), .ZN(n3197)
         );
  OAI22_X1 U1297 ( .A1(n419), .A2(n1583), .B1(n1737), .B2(n1804), .ZN(n3196)
         );
  OAI22_X1 U1298 ( .A1(n420), .A2(n1583), .B1(n1737), .B2(n1805), .ZN(n3195)
         );
  OAI22_X1 U1299 ( .A1(n421), .A2(n1583), .B1(n1737), .B2(n1806), .ZN(n3194)
         );
  OAI22_X1 U1300 ( .A1(n422), .A2(n1583), .B1(n1737), .B2(n1807), .ZN(n3193)
         );
  OAI22_X1 U1301 ( .A1(n423), .A2(n1583), .B1(n1737), .B2(n1808), .ZN(n3192)
         );
  OAI22_X1 U1302 ( .A1(n424), .A2(n1583), .B1(n1737), .B2(n1809), .ZN(n3191)
         );
  OAI22_X1 U1303 ( .A1(n425), .A2(n1583), .B1(n1737), .B2(n1810), .ZN(n3190)
         );
  OAI22_X1 U1304 ( .A1(n426), .A2(n1583), .B1(n1737), .B2(n1811), .ZN(n3189)
         );
  OAI22_X1 U1305 ( .A1(n427), .A2(n1583), .B1(n1737), .B2(n1812), .ZN(n3188)
         );
  OAI22_X1 U1306 ( .A1(n428), .A2(n1583), .B1(n1737), .B2(n1813), .ZN(n3187)
         );
  OAI22_X1 U1307 ( .A1(n429), .A2(n1583), .B1(n1666), .B2(n1814), .ZN(n3186)
         );
  OAI22_X1 U1308 ( .A1(n430), .A2(n1583), .B1(n1666), .B2(n1815), .ZN(n3185)
         );
  OAI22_X1 U1309 ( .A1(n431), .A2(n1583), .B1(n1666), .B2(n1816), .ZN(n3184)
         );
  OAI22_X1 U1310 ( .A1(n432), .A2(n1583), .B1(n1666), .B2(n1817), .ZN(n3183)
         );
  OAI22_X1 U1311 ( .A1(n433), .A2(n1583), .B1(n1666), .B2(n1818), .ZN(n3182)
         );
  OAI22_X1 U1312 ( .A1(n434), .A2(n1583), .B1(n1666), .B2(n1819), .ZN(n3181)
         );
  OAI22_X1 U1313 ( .A1(n435), .A2(n1583), .B1(n1666), .B2(n1820), .ZN(n3180)
         );
  OAI22_X1 U1314 ( .A1(n436), .A2(n1583), .B1(n1666), .B2(n1821), .ZN(n3179)
         );
  OAI22_X1 U1315 ( .A1(n437), .A2(n1583), .B1(n1666), .B2(n1822), .ZN(n3178)
         );
  OAI22_X1 U1316 ( .A1(n438), .A2(n1583), .B1(n1666), .B2(n1823), .ZN(n3177)
         );
  OAI22_X1 U1317 ( .A1(n439), .A2(n1583), .B1(n1666), .B2(n1824), .ZN(n3176)
         );
  OAI22_X1 U1318 ( .A1(n440), .A2(n1583), .B1(n1666), .B2(n1825), .ZN(n3175)
         );
  OAI22_X1 U1319 ( .A1(n441), .A2(n1738), .B1(n1666), .B2(n1826), .ZN(n3174)
         );
  OAI22_X1 U1320 ( .A1(n442), .A2(n1738), .B1(n1666), .B2(n1827), .ZN(n3173)
         );
  OAI22_X1 U1321 ( .A1(n443), .A2(n1583), .B1(n1666), .B2(n1828), .ZN(n3172)
         );
  OAI22_X1 U1322 ( .A1(n444), .A2(n1738), .B1(n1666), .B2(n1829), .ZN(n3171)
         );
  OAI22_X1 U1323 ( .A1(n445), .A2(n1738), .B1(n1737), .B2(n1830), .ZN(n3170)
         );
  OAI22_X1 U1324 ( .A1(n446), .A2(n1738), .B1(n1737), .B2(n1831), .ZN(n3169)
         );
  OAI22_X1 U1325 ( .A1(n447), .A2(n1738), .B1(n1737), .B2(n1832), .ZN(n3168)
         );
  OAI22_X1 U1326 ( .A1(n448), .A2(n1583), .B1(n1737), .B2(n1833), .ZN(n3167)
         );
  NAND2_X1 U1327 ( .A1(n1801), .A2(n1740), .ZN(n1739) );
  OAI22_X1 U1328 ( .A1(n449), .A2(n1603), .B1(n1741), .B2(n1802), .ZN(n3166)
         );
  OAI22_X1 U1329 ( .A1(n450), .A2(n1603), .B1(n1741), .B2(n1803), .ZN(n3165)
         );
  OAI22_X1 U1330 ( .A1(n451), .A2(n1603), .B1(n1741), .B2(n1804), .ZN(n3164)
         );
  OAI22_X1 U1331 ( .A1(n452), .A2(n1603), .B1(n1741), .B2(n1805), .ZN(n3163)
         );
  OAI22_X1 U1332 ( .A1(n453), .A2(n1603), .B1(n1741), .B2(n1806), .ZN(n3162)
         );
  OAI22_X1 U1333 ( .A1(n454), .A2(n1603), .B1(n1741), .B2(n1807), .ZN(n3161)
         );
  OAI22_X1 U1334 ( .A1(n455), .A2(n1603), .B1(n1741), .B2(n1808), .ZN(n3160)
         );
  OAI22_X1 U1335 ( .A1(n456), .A2(n1603), .B1(n1741), .B2(n1809), .ZN(n3159)
         );
  OAI22_X1 U1336 ( .A1(n457), .A2(n1603), .B1(n1741), .B2(n1810), .ZN(n3158)
         );
  OAI22_X1 U1337 ( .A1(n458), .A2(n1603), .B1(n1741), .B2(n1811), .ZN(n3157)
         );
  OAI22_X1 U1338 ( .A1(n459), .A2(n1603), .B1(n1741), .B2(n1812), .ZN(n3156)
         );
  OAI22_X1 U1339 ( .A1(n460), .A2(n1603), .B1(n1741), .B2(n1813), .ZN(n3155)
         );
  OAI22_X1 U1340 ( .A1(n461), .A2(n1603), .B1(n1667), .B2(n1814), .ZN(n3154)
         );
  OAI22_X1 U1341 ( .A1(n462), .A2(n1603), .B1(n1667), .B2(n1815), .ZN(n3153)
         );
  OAI22_X1 U1342 ( .A1(n463), .A2(n1603), .B1(n1667), .B2(n1816), .ZN(n3152)
         );
  OAI22_X1 U1343 ( .A1(n464), .A2(n1603), .B1(n1667), .B2(n1817), .ZN(n3151)
         );
  OAI22_X1 U1344 ( .A1(n465), .A2(n1603), .B1(n1667), .B2(n1818), .ZN(n3150)
         );
  OAI22_X1 U1345 ( .A1(n466), .A2(n1603), .B1(n1667), .B2(n1819), .ZN(n3149)
         );
  OAI22_X1 U1346 ( .A1(n467), .A2(n1603), .B1(n1667), .B2(n1820), .ZN(n3148)
         );
  OAI22_X1 U1347 ( .A1(n468), .A2(n1603), .B1(n1667), .B2(n1821), .ZN(n3147)
         );
  OAI22_X1 U1348 ( .A1(n469), .A2(n1603), .B1(n1667), .B2(n1822), .ZN(n3146)
         );
  OAI22_X1 U1349 ( .A1(n470), .A2(n1603), .B1(n1667), .B2(n1823), .ZN(n3145)
         );
  OAI22_X1 U1350 ( .A1(n471), .A2(n1603), .B1(n1667), .B2(n1824), .ZN(n3144)
         );
  OAI22_X1 U1351 ( .A1(n472), .A2(n1603), .B1(n1667), .B2(n1825), .ZN(n3143)
         );
  OAI22_X1 U1352 ( .A1(n473), .A2(n1742), .B1(n1667), .B2(n1826), .ZN(n3142)
         );
  OAI22_X1 U1353 ( .A1(n474), .A2(n1742), .B1(n1667), .B2(n1827), .ZN(n3141)
         );
  OAI22_X1 U1354 ( .A1(n475), .A2(n1603), .B1(n1667), .B2(n1828), .ZN(n3140)
         );
  OAI22_X1 U1355 ( .A1(n476), .A2(n1742), .B1(n1667), .B2(n1829), .ZN(n3139)
         );
  OAI22_X1 U1356 ( .A1(n477), .A2(n1742), .B1(n1741), .B2(n1830), .ZN(n3138)
         );
  OAI22_X1 U1357 ( .A1(n478), .A2(n1742), .B1(n1741), .B2(n1831), .ZN(n3137)
         );
  OAI22_X1 U1358 ( .A1(n479), .A2(n1742), .B1(n1741), .B2(n1832), .ZN(n3136)
         );
  OAI22_X1 U1359 ( .A1(n480), .A2(n1603), .B1(n1741), .B2(n1833), .ZN(n3135)
         );
  NAND2_X1 U1360 ( .A1(n1772), .A2(n1766), .ZN(n1744) );
  OAI22_X1 U1361 ( .A1(n481), .A2(n1602), .B1(n1745), .B2(n1802), .ZN(n3134)
         );
  OAI22_X1 U1362 ( .A1(n482), .A2(n1602), .B1(n1745), .B2(n1803), .ZN(n3133)
         );
  OAI22_X1 U1363 ( .A1(n483), .A2(n1602), .B1(n1745), .B2(n1804), .ZN(n3132)
         );
  OAI22_X1 U1364 ( .A1(n484), .A2(n1602), .B1(n1745), .B2(n1805), .ZN(n3131)
         );
  OAI22_X1 U1365 ( .A1(n485), .A2(n1602), .B1(n1745), .B2(n1806), .ZN(n3130)
         );
  OAI22_X1 U1366 ( .A1(n486), .A2(n1602), .B1(n1745), .B2(n1807), .ZN(n3129)
         );
  OAI22_X1 U1367 ( .A1(n487), .A2(n1602), .B1(n1745), .B2(n1808), .ZN(n3128)
         );
  OAI22_X1 U1368 ( .A1(n488), .A2(n1602), .B1(n1745), .B2(n1809), .ZN(n3127)
         );
  OAI22_X1 U1369 ( .A1(n489), .A2(n1602), .B1(n1745), .B2(n1810), .ZN(n3126)
         );
  OAI22_X1 U1370 ( .A1(n490), .A2(n1602), .B1(n1745), .B2(n1811), .ZN(n3125)
         );
  OAI22_X1 U1371 ( .A1(n491), .A2(n1602), .B1(n1745), .B2(n1812), .ZN(n3124)
         );
  OAI22_X1 U1372 ( .A1(n492), .A2(n1602), .B1(n1745), .B2(n1813), .ZN(n3123)
         );
  OAI22_X1 U1373 ( .A1(n493), .A2(n1602), .B1(n1745), .B2(n1814), .ZN(n3122)
         );
  OAI22_X1 U1374 ( .A1(n494), .A2(n1602), .B1(n1745), .B2(n1815), .ZN(n3121)
         );
  OAI22_X1 U1375 ( .A1(n495), .A2(n1602), .B1(n1745), .B2(n1816), .ZN(n3120)
         );
  OAI22_X1 U1376 ( .A1(n496), .A2(n1602), .B1(n1745), .B2(n1817), .ZN(n3119)
         );
  OAI22_X1 U1377 ( .A1(n497), .A2(n1602), .B1(n1745), .B2(n1818), .ZN(n3118)
         );
  OAI22_X1 U1378 ( .A1(n498), .A2(n1602), .B1(n1745), .B2(n1819), .ZN(n3117)
         );
  OAI22_X1 U1379 ( .A1(n499), .A2(n1602), .B1(n1745), .B2(n1820), .ZN(n3116)
         );
  OAI22_X1 U1380 ( .A1(n500), .A2(n1602), .B1(n1745), .B2(n1821), .ZN(n3115)
         );
  OAI22_X1 U1381 ( .A1(n501), .A2(n1602), .B1(n1745), .B2(n1822), .ZN(n3114)
         );
  OAI22_X1 U1382 ( .A1(n502), .A2(n1602), .B1(n1745), .B2(n1823), .ZN(n3113)
         );
  OAI22_X1 U1383 ( .A1(n503), .A2(n1602), .B1(n1745), .B2(n1824), .ZN(n3112)
         );
  OAI22_X1 U1384 ( .A1(n504), .A2(n1602), .B1(n1745), .B2(n1825), .ZN(n3111)
         );
  OAI22_X1 U1385 ( .A1(n505), .A2(n1746), .B1(n1745), .B2(n1826), .ZN(n3110)
         );
  OAI22_X1 U1386 ( .A1(n506), .A2(n1746), .B1(n1745), .B2(n1827), .ZN(n3109)
         );
  OAI22_X1 U1387 ( .A1(n507), .A2(n1602), .B1(n1745), .B2(n1828), .ZN(n3108)
         );
  OAI22_X1 U1388 ( .A1(n508), .A2(n1746), .B1(n1745), .B2(n1829), .ZN(n3107)
         );
  OAI22_X1 U1389 ( .A1(n509), .A2(n1746), .B1(n1745), .B2(n1830), .ZN(n3106)
         );
  OAI22_X1 U1390 ( .A1(n510), .A2(n1746), .B1(n1745), .B2(n1831), .ZN(n3105)
         );
  OAI22_X1 U1391 ( .A1(n511), .A2(n1746), .B1(n1745), .B2(n1832), .ZN(n3104)
         );
  OAI22_X1 U1392 ( .A1(n512), .A2(n1602), .B1(n1745), .B2(n1833), .ZN(n3103)
         );
  NAND2_X1 U1393 ( .A1(n1776), .A2(n1766), .ZN(n1747) );
  OAI22_X1 U1394 ( .A1(n513), .A2(n1610), .B1(n1748), .B2(n1802), .ZN(n3102)
         );
  OAI22_X1 U1395 ( .A1(n514), .A2(n1610), .B1(n1748), .B2(n1803), .ZN(n3101)
         );
  OAI22_X1 U1396 ( .A1(n515), .A2(n1610), .B1(n1748), .B2(n1804), .ZN(n3100)
         );
  OAI22_X1 U1397 ( .A1(n516), .A2(n1610), .B1(n1748), .B2(n1805), .ZN(n3099)
         );
  OAI22_X1 U1398 ( .A1(n517), .A2(n1610), .B1(n1748), .B2(n1806), .ZN(n3098)
         );
  OAI22_X1 U1399 ( .A1(n518), .A2(n1610), .B1(n1748), .B2(n1807), .ZN(n3097)
         );
  OAI22_X1 U1400 ( .A1(n519), .A2(n1610), .B1(n1748), .B2(n1808), .ZN(n3096)
         );
  OAI22_X1 U1401 ( .A1(n520), .A2(n1610), .B1(n1748), .B2(n1809), .ZN(n3095)
         );
  OAI22_X1 U1402 ( .A1(n521), .A2(n1610), .B1(n1748), .B2(n1810), .ZN(n3094)
         );
  OAI22_X1 U1403 ( .A1(n522), .A2(n1610), .B1(n1748), .B2(n1811), .ZN(n3093)
         );
  OAI22_X1 U1404 ( .A1(n523), .A2(n1610), .B1(n1748), .B2(n1812), .ZN(n3092)
         );
  OAI22_X1 U1405 ( .A1(n524), .A2(n1610), .B1(n1748), .B2(n1813), .ZN(n3091)
         );
  OAI22_X1 U1406 ( .A1(n525), .A2(n1610), .B1(n1668), .B2(n1814), .ZN(n3090)
         );
  OAI22_X1 U1407 ( .A1(n526), .A2(n1610), .B1(n1668), .B2(n1815), .ZN(n3089)
         );
  OAI22_X1 U1408 ( .A1(n527), .A2(n1610), .B1(n1668), .B2(n1816), .ZN(n3088)
         );
  OAI22_X1 U1409 ( .A1(n528), .A2(n1610), .B1(n1668), .B2(n1817), .ZN(n3087)
         );
  OAI22_X1 U1410 ( .A1(n529), .A2(n1610), .B1(n1668), .B2(n1818), .ZN(n3086)
         );
  OAI22_X1 U1411 ( .A1(n530), .A2(n1610), .B1(n1668), .B2(n1819), .ZN(n3085)
         );
  OAI22_X1 U1412 ( .A1(n531), .A2(n1610), .B1(n1668), .B2(n1820), .ZN(n3084)
         );
  OAI22_X1 U1413 ( .A1(n532), .A2(n1610), .B1(n1668), .B2(n1821), .ZN(n3083)
         );
  OAI22_X1 U1414 ( .A1(n533), .A2(n1610), .B1(n1668), .B2(n1822), .ZN(n3082)
         );
  OAI22_X1 U1415 ( .A1(n534), .A2(n1610), .B1(n1668), .B2(n1823), .ZN(n3081)
         );
  OAI22_X1 U1416 ( .A1(n535), .A2(n1610), .B1(n1668), .B2(n1824), .ZN(n3080)
         );
  OAI22_X1 U1417 ( .A1(n536), .A2(n1610), .B1(n1668), .B2(n1825), .ZN(n3079)
         );
  OAI22_X1 U1418 ( .A1(n537), .A2(n1749), .B1(n1668), .B2(n1826), .ZN(n3078)
         );
  OAI22_X1 U1419 ( .A1(n538), .A2(n1749), .B1(n1748), .B2(n1827), .ZN(n3077)
         );
  OAI22_X1 U1420 ( .A1(n539), .A2(n1610), .B1(n1668), .B2(n1828), .ZN(n3076)
         );
  OAI22_X1 U1421 ( .A1(n540), .A2(n1749), .B1(n1668), .B2(n1829), .ZN(n3075)
         );
  OAI22_X1 U1422 ( .A1(n541), .A2(n1749), .B1(n1748), .B2(n1830), .ZN(n3074)
         );
  OAI22_X1 U1423 ( .A1(n542), .A2(n1749), .B1(n1748), .B2(n1831), .ZN(n3073)
         );
  OAI22_X1 U1424 ( .A1(n543), .A2(n1749), .B1(n1668), .B2(n1832), .ZN(n3072)
         );
  OAI22_X1 U1425 ( .A1(n544), .A2(n1610), .B1(n1668), .B2(n1833), .ZN(n3071)
         );
  NAND2_X1 U1426 ( .A1(n1780), .A2(n1766), .ZN(n1750) );
  NAND3_X1 U1427 ( .A1(rst), .A2(n1780), .A3(n1766), .ZN(n1751) );
  OAI22_X1 U1428 ( .A1(n545), .A2(n1585), .B1(n1619), .B2(n1802), .ZN(n3070)
         );
  OAI22_X1 U1429 ( .A1(n546), .A2(n1585), .B1(n1619), .B2(n1803), .ZN(n3069)
         );
  OAI22_X1 U1430 ( .A1(n547), .A2(n1585), .B1(n1619), .B2(n1804), .ZN(n3068)
         );
  OAI22_X1 U1431 ( .A1(n548), .A2(n1585), .B1(n1619), .B2(n1805), .ZN(n3067)
         );
  OAI22_X1 U1432 ( .A1(n549), .A2(n1585), .B1(n1619), .B2(n1806), .ZN(n3066)
         );
  OAI22_X1 U1433 ( .A1(n550), .A2(n1585), .B1(n1619), .B2(n1807), .ZN(n3065)
         );
  OAI22_X1 U1434 ( .A1(n551), .A2(n1585), .B1(n1619), .B2(n1808), .ZN(n3064)
         );
  OAI22_X1 U1435 ( .A1(n552), .A2(n1585), .B1(n1619), .B2(n1809), .ZN(n3063)
         );
  OAI22_X1 U1436 ( .A1(n553), .A2(n1585), .B1(n1619), .B2(n1810), .ZN(n3062)
         );
  OAI22_X1 U1437 ( .A1(n554), .A2(n1585), .B1(n1619), .B2(n1811), .ZN(n3061)
         );
  OAI22_X1 U1438 ( .A1(n555), .A2(n1585), .B1(n1619), .B2(n1812), .ZN(n3060)
         );
  OAI22_X1 U1439 ( .A1(n556), .A2(n1585), .B1(n1619), .B2(n1813), .ZN(n3059)
         );
  OAI22_X1 U1440 ( .A1(n557), .A2(n1585), .B1(n1619), .B2(n1814), .ZN(n3058)
         );
  OAI22_X1 U1441 ( .A1(n558), .A2(n1585), .B1(n1619), .B2(n1815), .ZN(n3057)
         );
  OAI22_X1 U1442 ( .A1(n559), .A2(n1585), .B1(n1619), .B2(n1816), .ZN(n3056)
         );
  OAI22_X1 U1443 ( .A1(n560), .A2(n1585), .B1(n1619), .B2(n1817), .ZN(n3055)
         );
  OAI22_X1 U1444 ( .A1(n561), .A2(n1585), .B1(n1619), .B2(n1818), .ZN(n3054)
         );
  OAI22_X1 U1445 ( .A1(n562), .A2(n1585), .B1(n1619), .B2(n1819), .ZN(n3053)
         );
  OAI22_X1 U1446 ( .A1(n563), .A2(n1585), .B1(n1619), .B2(n1820), .ZN(n3052)
         );
  OAI22_X1 U1447 ( .A1(n564), .A2(n1585), .B1(n1619), .B2(n1821), .ZN(n3051)
         );
  OAI22_X1 U1448 ( .A1(n565), .A2(n1585), .B1(n1619), .B2(n1822), .ZN(n3050)
         );
  OAI22_X1 U1449 ( .A1(n566), .A2(n1585), .B1(n1619), .B2(n1823), .ZN(n3049)
         );
  OAI22_X1 U1450 ( .A1(n567), .A2(n1585), .B1(n1619), .B2(n1824), .ZN(n3048)
         );
  OAI22_X1 U1451 ( .A1(n568), .A2(n1585), .B1(n1619), .B2(n1825), .ZN(n3047)
         );
  OAI22_X1 U1452 ( .A1(n569), .A2(n1752), .B1(n1619), .B2(n1826), .ZN(n3046)
         );
  OAI22_X1 U1453 ( .A1(n570), .A2(n1752), .B1(n1619), .B2(n1827), .ZN(n3045)
         );
  OAI22_X1 U1454 ( .A1(n571), .A2(n1585), .B1(n1619), .B2(n1828), .ZN(n3044)
         );
  OAI22_X1 U1455 ( .A1(n572), .A2(n1752), .B1(n1619), .B2(n1829), .ZN(n3043)
         );
  OAI22_X1 U1456 ( .A1(n573), .A2(n1752), .B1(n1751), .B2(n1830), .ZN(n3042)
         );
  OAI22_X1 U1457 ( .A1(n574), .A2(n1752), .B1(n1751), .B2(n1831), .ZN(n3041)
         );
  OAI22_X1 U1458 ( .A1(n575), .A2(n1752), .B1(n1751), .B2(n1832), .ZN(n3040)
         );
  OAI22_X1 U1459 ( .A1(n576), .A2(n1585), .B1(n1751), .B2(n1833), .ZN(n3039)
         );
  NAND2_X1 U1460 ( .A1(n1784), .A2(n1766), .ZN(n1753) );
  OAI22_X1 U1461 ( .A1(n577), .A2(n1607), .B1(n1754), .B2(n1802), .ZN(n3038)
         );
  OAI22_X1 U1462 ( .A1(n578), .A2(n1607), .B1(n1754), .B2(n1803), .ZN(n3037)
         );
  OAI22_X1 U1463 ( .A1(n579), .A2(n1607), .B1(n1754), .B2(n1804), .ZN(n3036)
         );
  OAI22_X1 U1464 ( .A1(n580), .A2(n1607), .B1(n1754), .B2(n1805), .ZN(n3035)
         );
  OAI22_X1 U1465 ( .A1(n581), .A2(n1607), .B1(n1754), .B2(n1806), .ZN(n3034)
         );
  OAI22_X1 U1466 ( .A1(n582), .A2(n1607), .B1(n1754), .B2(n1807), .ZN(n3033)
         );
  OAI22_X1 U1467 ( .A1(n583), .A2(n1607), .B1(n1754), .B2(n1808), .ZN(n3032)
         );
  OAI22_X1 U1468 ( .A1(n584), .A2(n1607), .B1(n1754), .B2(n1809), .ZN(n3031)
         );
  OAI22_X1 U1469 ( .A1(n585), .A2(n1607), .B1(n1754), .B2(n1810), .ZN(n3030)
         );
  OAI22_X1 U1470 ( .A1(n586), .A2(n1607), .B1(n1754), .B2(n1811), .ZN(n3029)
         );
  OAI22_X1 U1471 ( .A1(n587), .A2(n1607), .B1(n1754), .B2(n1812), .ZN(n3028)
         );
  OAI22_X1 U1472 ( .A1(n588), .A2(n1607), .B1(n1754), .B2(n1813), .ZN(n3027)
         );
  OAI22_X1 U1473 ( .A1(n589), .A2(n1607), .B1(n1669), .B2(n1814), .ZN(n3026)
         );
  OAI22_X1 U1474 ( .A1(n590), .A2(n1607), .B1(n1669), .B2(n1815), .ZN(n3025)
         );
  OAI22_X1 U1475 ( .A1(n591), .A2(n1607), .B1(n1669), .B2(n1816), .ZN(n3024)
         );
  OAI22_X1 U1476 ( .A1(n592), .A2(n1607), .B1(n1669), .B2(n1817), .ZN(n3023)
         );
  OAI22_X1 U1477 ( .A1(n593), .A2(n1607), .B1(n1669), .B2(n1818), .ZN(n3022)
         );
  OAI22_X1 U1478 ( .A1(n594), .A2(n1607), .B1(n1669), .B2(n1819), .ZN(n3021)
         );
  OAI22_X1 U1479 ( .A1(n595), .A2(n1607), .B1(n1669), .B2(n1820), .ZN(n3020)
         );
  OAI22_X1 U1480 ( .A1(n596), .A2(n1607), .B1(n1669), .B2(n1821), .ZN(n3019)
         );
  OAI22_X1 U1481 ( .A1(n597), .A2(n1607), .B1(n1669), .B2(n1822), .ZN(n3018)
         );
  OAI22_X1 U1482 ( .A1(n598), .A2(n1607), .B1(n1669), .B2(n1823), .ZN(n3017)
         );
  OAI22_X1 U1483 ( .A1(n599), .A2(n1607), .B1(n1669), .B2(n1824), .ZN(n3016)
         );
  OAI22_X1 U1484 ( .A1(n600), .A2(n1607), .B1(n1669), .B2(n1825), .ZN(n3015)
         );
  OAI22_X1 U1485 ( .A1(n601), .A2(n1755), .B1(n1669), .B2(n1826), .ZN(n3014)
         );
  OAI22_X1 U1486 ( .A1(n602), .A2(n1755), .B1(n1754), .B2(n1827), .ZN(n3013)
         );
  OAI22_X1 U1487 ( .A1(n603), .A2(n1607), .B1(n1669), .B2(n1828), .ZN(n3012)
         );
  OAI22_X1 U1488 ( .A1(n604), .A2(n1755), .B1(n1669), .B2(n1829), .ZN(n3011)
         );
  OAI22_X1 U1489 ( .A1(n605), .A2(n1755), .B1(n1754), .B2(n1830), .ZN(n3010)
         );
  OAI22_X1 U1490 ( .A1(n606), .A2(n1755), .B1(n1754), .B2(n1831), .ZN(n3009)
         );
  OAI22_X1 U1491 ( .A1(n607), .A2(n1755), .B1(n1754), .B2(n1832), .ZN(n3008)
         );
  OAI22_X1 U1492 ( .A1(n608), .A2(n1607), .B1(n1754), .B2(n1833), .ZN(n3007)
         );
  NAND2_X1 U1493 ( .A1(n1788), .A2(n1766), .ZN(n1756) );
  OAI22_X1 U1494 ( .A1(n609), .A2(n1608), .B1(n1757), .B2(n1802), .ZN(n3006)
         );
  OAI22_X1 U1495 ( .A1(n610), .A2(n1608), .B1(n1757), .B2(n1803), .ZN(n3005)
         );
  OAI22_X1 U1496 ( .A1(n611), .A2(n1608), .B1(n1757), .B2(n1804), .ZN(n3004)
         );
  OAI22_X1 U1497 ( .A1(n612), .A2(n1608), .B1(n1757), .B2(n1805), .ZN(n3003)
         );
  OAI22_X1 U1498 ( .A1(n613), .A2(n1608), .B1(n1757), .B2(n1806), .ZN(n3002)
         );
  OAI22_X1 U1499 ( .A1(n614), .A2(n1608), .B1(n1757), .B2(n1807), .ZN(n3001)
         );
  OAI22_X1 U1500 ( .A1(n615), .A2(n1608), .B1(n1757), .B2(n1808), .ZN(n3000)
         );
  OAI22_X1 U1501 ( .A1(n616), .A2(n1608), .B1(n1757), .B2(n1809), .ZN(n2999)
         );
  OAI22_X1 U1502 ( .A1(n617), .A2(n1608), .B1(n1757), .B2(n1810), .ZN(n2998)
         );
  OAI22_X1 U1503 ( .A1(n618), .A2(n1608), .B1(n1757), .B2(n1811), .ZN(n2997)
         );
  OAI22_X1 U1504 ( .A1(n619), .A2(n1608), .B1(n1757), .B2(n1812), .ZN(n2996)
         );
  OAI22_X1 U1505 ( .A1(n620), .A2(n1608), .B1(n1757), .B2(n1813), .ZN(n2995)
         );
  OAI22_X1 U1506 ( .A1(n621), .A2(n1608), .B1(n1670), .B2(n1814), .ZN(n2994)
         );
  OAI22_X1 U1507 ( .A1(n622), .A2(n1608), .B1(n1670), .B2(n1815), .ZN(n2993)
         );
  OAI22_X1 U1508 ( .A1(n623), .A2(n1608), .B1(n1670), .B2(n1816), .ZN(n2992)
         );
  OAI22_X1 U1509 ( .A1(n624), .A2(n1608), .B1(n1670), .B2(n1817), .ZN(n2991)
         );
  OAI22_X1 U1510 ( .A1(n625), .A2(n1608), .B1(n1670), .B2(n1818), .ZN(n2990)
         );
  OAI22_X1 U1511 ( .A1(n626), .A2(n1608), .B1(n1670), .B2(n1819), .ZN(n2989)
         );
  OAI22_X1 U1512 ( .A1(n627), .A2(n1608), .B1(n1670), .B2(n1820), .ZN(n2988)
         );
  OAI22_X1 U1513 ( .A1(n628), .A2(n1608), .B1(n1670), .B2(n1821), .ZN(n2987)
         );
  OAI22_X1 U1514 ( .A1(n629), .A2(n1608), .B1(n1670), .B2(n1822), .ZN(n2986)
         );
  OAI22_X1 U1515 ( .A1(n630), .A2(n1608), .B1(n1670), .B2(n1823), .ZN(n2985)
         );
  OAI22_X1 U1516 ( .A1(n631), .A2(n1608), .B1(n1670), .B2(n1824), .ZN(n2984)
         );
  OAI22_X1 U1517 ( .A1(n632), .A2(n1608), .B1(n1670), .B2(n1825), .ZN(n2983)
         );
  OAI22_X1 U1518 ( .A1(n633), .A2(n1758), .B1(n1670), .B2(n1826), .ZN(n2982)
         );
  OAI22_X1 U1519 ( .A1(n634), .A2(n1758), .B1(n1757), .B2(n1827), .ZN(n2981)
         );
  OAI22_X1 U1520 ( .A1(n635), .A2(n1608), .B1(n1670), .B2(n1828), .ZN(n2980)
         );
  OAI22_X1 U1521 ( .A1(n636), .A2(n1758), .B1(n1670), .B2(n1829), .ZN(n2979)
         );
  OAI22_X1 U1522 ( .A1(n637), .A2(n1758), .B1(n1757), .B2(n1830), .ZN(n2978)
         );
  OAI22_X1 U1523 ( .A1(n638), .A2(n1758), .B1(n1757), .B2(n1831), .ZN(n2977)
         );
  OAI22_X1 U1524 ( .A1(n639), .A2(n1758), .B1(n1670), .B2(n1832), .ZN(n2976)
         );
  OAI22_X1 U1525 ( .A1(n640), .A2(n1608), .B1(n1670), .B2(n1833), .ZN(n2975)
         );
  NAND2_X1 U1526 ( .A1(n1792), .A2(n1766), .ZN(n1759) );
  OAI22_X1 U1527 ( .A1(n641), .A2(n1613), .B1(n1760), .B2(n1802), .ZN(n2974)
         );
  OAI22_X1 U1528 ( .A1(n642), .A2(n1613), .B1(n1760), .B2(n1803), .ZN(n2973)
         );
  OAI22_X1 U1529 ( .A1(n643), .A2(n1613), .B1(n1760), .B2(n1804), .ZN(n2972)
         );
  OAI22_X1 U1530 ( .A1(n644), .A2(n1613), .B1(n1760), .B2(n1805), .ZN(n2971)
         );
  OAI22_X1 U1531 ( .A1(n645), .A2(n1613), .B1(n1760), .B2(n1806), .ZN(n2970)
         );
  OAI22_X1 U1532 ( .A1(n646), .A2(n1613), .B1(n1760), .B2(n1807), .ZN(n2969)
         );
  OAI22_X1 U1533 ( .A1(n647), .A2(n1613), .B1(n1760), .B2(n1808), .ZN(n2968)
         );
  OAI22_X1 U1534 ( .A1(n648), .A2(n1613), .B1(n1760), .B2(n1809), .ZN(n2967)
         );
  OAI22_X1 U1535 ( .A1(n649), .A2(n1613), .B1(n1760), .B2(n1810), .ZN(n2966)
         );
  OAI22_X1 U1536 ( .A1(n650), .A2(n1613), .B1(n1760), .B2(n1811), .ZN(n2965)
         );
  OAI22_X1 U1537 ( .A1(n651), .A2(n1613), .B1(n1760), .B2(n1812), .ZN(n2964)
         );
  OAI22_X1 U1538 ( .A1(n652), .A2(n1613), .B1(n1760), .B2(n1813), .ZN(n2963)
         );
  OAI22_X1 U1539 ( .A1(n653), .A2(n1613), .B1(n1671), .B2(n1814), .ZN(n2962)
         );
  OAI22_X1 U1540 ( .A1(n654), .A2(n1613), .B1(n1671), .B2(n1815), .ZN(n2961)
         );
  OAI22_X1 U1541 ( .A1(n655), .A2(n1613), .B1(n1671), .B2(n1816), .ZN(n2960)
         );
  OAI22_X1 U1542 ( .A1(n656), .A2(n1613), .B1(n1671), .B2(n1817), .ZN(n2959)
         );
  OAI22_X1 U1543 ( .A1(n657), .A2(n1613), .B1(n1671), .B2(n1818), .ZN(n2958)
         );
  OAI22_X1 U1544 ( .A1(n658), .A2(n1613), .B1(n1671), .B2(n1819), .ZN(n2957)
         );
  OAI22_X1 U1545 ( .A1(n659), .A2(n1613), .B1(n1671), .B2(n1820), .ZN(n2956)
         );
  OAI22_X1 U1546 ( .A1(n660), .A2(n1613), .B1(n1671), .B2(n1821), .ZN(n2955)
         );
  OAI22_X1 U1547 ( .A1(n661), .A2(n1613), .B1(n1671), .B2(n1822), .ZN(n2954)
         );
  OAI22_X1 U1548 ( .A1(n662), .A2(n1613), .B1(n1671), .B2(n1823), .ZN(n2953)
         );
  OAI22_X1 U1549 ( .A1(n663), .A2(n1613), .B1(n1671), .B2(n1824), .ZN(n2952)
         );
  OAI22_X1 U1550 ( .A1(n664), .A2(n1613), .B1(n1671), .B2(n1825), .ZN(n2951)
         );
  OAI22_X1 U1551 ( .A1(n665), .A2(n1761), .B1(n1671), .B2(n1826), .ZN(n2950)
         );
  OAI22_X1 U1552 ( .A1(n666), .A2(n1761), .B1(n1760), .B2(n1827), .ZN(n2949)
         );
  OAI22_X1 U1553 ( .A1(n667), .A2(n1613), .B1(n1671), .B2(n1828), .ZN(n2948)
         );
  OAI22_X1 U1554 ( .A1(n668), .A2(n1761), .B1(n1671), .B2(n1829), .ZN(n2947)
         );
  OAI22_X1 U1555 ( .A1(n669), .A2(n1761), .B1(n1760), .B2(n1830), .ZN(n2946)
         );
  OAI22_X1 U1556 ( .A1(n670), .A2(n1761), .B1(n1760), .B2(n1831), .ZN(n2945)
         );
  OAI22_X1 U1557 ( .A1(n671), .A2(n1761), .B1(n1671), .B2(n1832), .ZN(n2944)
         );
  OAI22_X1 U1558 ( .A1(n672), .A2(n1613), .B1(n1671), .B2(n1833), .ZN(n2943)
         );
  NAND2_X1 U1559 ( .A1(n1796), .A2(n1766), .ZN(n1762) );
  NAND3_X1 U1560 ( .A1(rst), .A2(n1796), .A3(n1766), .ZN(n1763) );
  OAI22_X1 U1561 ( .A1(n673), .A2(n1591), .B1(n1618), .B2(n1802), .ZN(n2942)
         );
  OAI22_X1 U1562 ( .A1(n674), .A2(n1591), .B1(n1618), .B2(n1803), .ZN(n2941)
         );
  OAI22_X1 U1563 ( .A1(n675), .A2(n1591), .B1(n1618), .B2(n1804), .ZN(n2940)
         );
  OAI22_X1 U1564 ( .A1(n676), .A2(n1591), .B1(n1618), .B2(n1805), .ZN(n2939)
         );
  OAI22_X1 U1565 ( .A1(n677), .A2(n1591), .B1(n1618), .B2(n1806), .ZN(n2938)
         );
  OAI22_X1 U1566 ( .A1(n678), .A2(n1591), .B1(n1618), .B2(n1807), .ZN(n2937)
         );
  OAI22_X1 U1567 ( .A1(n679), .A2(n1591), .B1(n1618), .B2(n1808), .ZN(n2936)
         );
  OAI22_X1 U1568 ( .A1(n680), .A2(n1591), .B1(n1618), .B2(n1809), .ZN(n2935)
         );
  OAI22_X1 U1569 ( .A1(n681), .A2(n1591), .B1(n1618), .B2(n1810), .ZN(n2934)
         );
  OAI22_X1 U1570 ( .A1(n682), .A2(n1591), .B1(n1618), .B2(n1811), .ZN(n2933)
         );
  OAI22_X1 U1571 ( .A1(n683), .A2(n1591), .B1(n1618), .B2(n1812), .ZN(n2932)
         );
  OAI22_X1 U1572 ( .A1(n684), .A2(n1591), .B1(n1618), .B2(n1813), .ZN(n2931)
         );
  OAI22_X1 U1573 ( .A1(n685), .A2(n1591), .B1(n1618), .B2(n1814), .ZN(n2930)
         );
  OAI22_X1 U1574 ( .A1(n686), .A2(n1591), .B1(n1618), .B2(n1815), .ZN(n2929)
         );
  OAI22_X1 U1575 ( .A1(n687), .A2(n1591), .B1(n1618), .B2(n1816), .ZN(n2928)
         );
  OAI22_X1 U1576 ( .A1(n688), .A2(n1591), .B1(n1618), .B2(n1817), .ZN(n2927)
         );
  OAI22_X1 U1577 ( .A1(n689), .A2(n1591), .B1(n1618), .B2(n1818), .ZN(n2926)
         );
  OAI22_X1 U1578 ( .A1(n690), .A2(n1591), .B1(n1618), .B2(n1819), .ZN(n2925)
         );
  OAI22_X1 U1579 ( .A1(n691), .A2(n1591), .B1(n1618), .B2(n1820), .ZN(n2924)
         );
  OAI22_X1 U1580 ( .A1(n692), .A2(n1591), .B1(n1618), .B2(n1821), .ZN(n2923)
         );
  OAI22_X1 U1581 ( .A1(n693), .A2(n1591), .B1(n1618), .B2(n1822), .ZN(n2922)
         );
  OAI22_X1 U1582 ( .A1(n694), .A2(n1591), .B1(n1618), .B2(n1823), .ZN(n2921)
         );
  OAI22_X1 U1583 ( .A1(n695), .A2(n1591), .B1(n1618), .B2(n1824), .ZN(n2920)
         );
  OAI22_X1 U1584 ( .A1(n696), .A2(n1591), .B1(n1618), .B2(n1825), .ZN(n2919)
         );
  OAI22_X1 U1585 ( .A1(n697), .A2(n1764), .B1(n1618), .B2(n1826), .ZN(n2918)
         );
  OAI22_X1 U1586 ( .A1(n698), .A2(n1764), .B1(n1618), .B2(n1827), .ZN(n2917)
         );
  OAI22_X1 U1587 ( .A1(n699), .A2(n1591), .B1(n1618), .B2(n1828), .ZN(n2916)
         );
  OAI22_X1 U1588 ( .A1(n700), .A2(n1764), .B1(n1618), .B2(n1829), .ZN(n2915)
         );
  OAI22_X1 U1589 ( .A1(n701), .A2(n1764), .B1(n1763), .B2(n1830), .ZN(n2914)
         );
  OAI22_X1 U1590 ( .A1(n702), .A2(n1764), .B1(n1763), .B2(n1831), .ZN(n2913)
         );
  OAI22_X1 U1591 ( .A1(n703), .A2(n1764), .B1(n1763), .B2(n1832), .ZN(n2912)
         );
  OAI22_X1 U1592 ( .A1(n704), .A2(n1591), .B1(n1763), .B2(n1833), .ZN(n2911)
         );
  NAND2_X1 U1593 ( .A1(n1801), .A2(n1766), .ZN(n1765) );
  OAI22_X1 U1594 ( .A1(n705), .A2(n1605), .B1(n1767), .B2(n1802), .ZN(n2910)
         );
  OAI22_X1 U1595 ( .A1(n706), .A2(n1605), .B1(n1767), .B2(n1803), .ZN(n2909)
         );
  OAI22_X1 U1596 ( .A1(n707), .A2(n1605), .B1(n1767), .B2(n1804), .ZN(n2908)
         );
  OAI22_X1 U1597 ( .A1(n708), .A2(n1605), .B1(n1767), .B2(n1805), .ZN(n2907)
         );
  OAI22_X1 U1598 ( .A1(n709), .A2(n1605), .B1(n1767), .B2(n1806), .ZN(n2906)
         );
  OAI22_X1 U1599 ( .A1(n710), .A2(n1605), .B1(n1767), .B2(n1807), .ZN(n2905)
         );
  OAI22_X1 U1600 ( .A1(n711), .A2(n1605), .B1(n1767), .B2(n1808), .ZN(n2904)
         );
  OAI22_X1 U1601 ( .A1(n712), .A2(n1605), .B1(n1767), .B2(n1809), .ZN(n2903)
         );
  OAI22_X1 U1602 ( .A1(n713), .A2(n1605), .B1(n1767), .B2(n1810), .ZN(n2902)
         );
  OAI22_X1 U1603 ( .A1(n714), .A2(n1605), .B1(n1767), .B2(n1811), .ZN(n2901)
         );
  OAI22_X1 U1604 ( .A1(n715), .A2(n1605), .B1(n1767), .B2(n1812), .ZN(n2900)
         );
  OAI22_X1 U1605 ( .A1(n716), .A2(n1605), .B1(n1767), .B2(n1813), .ZN(n2899)
         );
  OAI22_X1 U1606 ( .A1(n717), .A2(n1605), .B1(n1672), .B2(n1814), .ZN(n2898)
         );
  OAI22_X1 U1607 ( .A1(n718), .A2(n1605), .B1(n1672), .B2(n1815), .ZN(n2897)
         );
  OAI22_X1 U1608 ( .A1(n719), .A2(n1605), .B1(n1672), .B2(n1816), .ZN(n2896)
         );
  OAI22_X1 U1609 ( .A1(n720), .A2(n1605), .B1(n1672), .B2(n1817), .ZN(n2895)
         );
  OAI22_X1 U1610 ( .A1(n721), .A2(n1605), .B1(n1672), .B2(n1818), .ZN(n2894)
         );
  OAI22_X1 U1611 ( .A1(n722), .A2(n1605), .B1(n1672), .B2(n1819), .ZN(n2893)
         );
  OAI22_X1 U1612 ( .A1(n723), .A2(n1605), .B1(n1672), .B2(n1820), .ZN(n2892)
         );
  OAI22_X1 U1613 ( .A1(n724), .A2(n1605), .B1(n1672), .B2(n1821), .ZN(n2891)
         );
  OAI22_X1 U1614 ( .A1(n725), .A2(n1605), .B1(n1672), .B2(n1822), .ZN(n2890)
         );
  OAI22_X1 U1615 ( .A1(n726), .A2(n1605), .B1(n1672), .B2(n1823), .ZN(n2889)
         );
  OAI22_X1 U1616 ( .A1(n727), .A2(n1605), .B1(n1672), .B2(n1824), .ZN(n2888)
         );
  OAI22_X1 U1617 ( .A1(n728), .A2(n1605), .B1(n1672), .B2(n1825), .ZN(n2887)
         );
  OAI22_X1 U1618 ( .A1(n729), .A2(n1768), .B1(n1672), .B2(n1826), .ZN(n2886)
         );
  OAI22_X1 U1619 ( .A1(n730), .A2(n1768), .B1(n1767), .B2(n1827), .ZN(n2885)
         );
  OAI22_X1 U1620 ( .A1(n731), .A2(n1605), .B1(n1672), .B2(n1828), .ZN(n2884)
         );
  OAI22_X1 U1621 ( .A1(n732), .A2(n1768), .B1(n1672), .B2(n1829), .ZN(n2883)
         );
  OAI22_X1 U1622 ( .A1(n733), .A2(n1768), .B1(n1767), .B2(n1830), .ZN(n2882)
         );
  OAI22_X1 U1623 ( .A1(n734), .A2(n1768), .B1(n1767), .B2(n1831), .ZN(n2881)
         );
  OAI22_X1 U1624 ( .A1(n735), .A2(n1768), .B1(n1767), .B2(n1832), .ZN(n2880)
         );
  OAI22_X1 U1625 ( .A1(n736), .A2(n1605), .B1(n1767), .B2(n1833), .ZN(n2879)
         );
  NAND2_X1 U1626 ( .A1(n1772), .A2(n1800), .ZN(n1771) );
  OAI22_X1 U1627 ( .A1(n737), .A2(n1612), .B1(n1773), .B2(n1802), .ZN(n2878)
         );
  OAI22_X1 U1628 ( .A1(n738), .A2(n1612), .B1(n1773), .B2(n1803), .ZN(n2877)
         );
  OAI22_X1 U1629 ( .A1(n739), .A2(n1612), .B1(n1773), .B2(n1804), .ZN(n2876)
         );
  OAI22_X1 U1630 ( .A1(n740), .A2(n1612), .B1(n1773), .B2(n1805), .ZN(n2875)
         );
  OAI22_X1 U1631 ( .A1(n741), .A2(n1612), .B1(n1773), .B2(n1806), .ZN(n2874)
         );
  OAI22_X1 U1632 ( .A1(n742), .A2(n1612), .B1(n1773), .B2(n1807), .ZN(n2873)
         );
  OAI22_X1 U1633 ( .A1(n743), .A2(n1612), .B1(n1773), .B2(n1808), .ZN(n2872)
         );
  OAI22_X1 U1634 ( .A1(n744), .A2(n1612), .B1(n1773), .B2(n1809), .ZN(n2871)
         );
  OAI22_X1 U1635 ( .A1(n745), .A2(n1612), .B1(n1773), .B2(n1810), .ZN(n2870)
         );
  OAI22_X1 U1636 ( .A1(n746), .A2(n1612), .B1(n1773), .B2(n1811), .ZN(n2869)
         );
  OAI22_X1 U1637 ( .A1(n747), .A2(n1612), .B1(n1773), .B2(n1812), .ZN(n2868)
         );
  OAI22_X1 U1638 ( .A1(n748), .A2(n1612), .B1(n1773), .B2(n1813), .ZN(n2867)
         );
  OAI22_X1 U1639 ( .A1(n749), .A2(n1612), .B1(n1673), .B2(n1814), .ZN(n2866)
         );
  OAI22_X1 U1640 ( .A1(n750), .A2(n1612), .B1(n1673), .B2(n1815), .ZN(n2865)
         );
  OAI22_X1 U1641 ( .A1(n751), .A2(n1612), .B1(n1673), .B2(n1816), .ZN(n2864)
         );
  OAI22_X1 U1642 ( .A1(n752), .A2(n1612), .B1(n1673), .B2(n1817), .ZN(n2863)
         );
  OAI22_X1 U1643 ( .A1(n753), .A2(n1612), .B1(n1673), .B2(n1818), .ZN(n2862)
         );
  OAI22_X1 U1644 ( .A1(n754), .A2(n1612), .B1(n1673), .B2(n1819), .ZN(n2861)
         );
  OAI22_X1 U1645 ( .A1(n755), .A2(n1612), .B1(n1673), .B2(n1820), .ZN(n2860)
         );
  OAI22_X1 U1646 ( .A1(n756), .A2(n1612), .B1(n1673), .B2(n1821), .ZN(n2859)
         );
  OAI22_X1 U1647 ( .A1(n757), .A2(n1612), .B1(n1673), .B2(n1822), .ZN(n2858)
         );
  OAI22_X1 U1648 ( .A1(n758), .A2(n1612), .B1(n1673), .B2(n1823), .ZN(n2857)
         );
  OAI22_X1 U1649 ( .A1(n759), .A2(n1612), .B1(n1673), .B2(n1824), .ZN(n2856)
         );
  OAI22_X1 U1650 ( .A1(n760), .A2(n1612), .B1(n1673), .B2(n1825), .ZN(n2855)
         );
  OAI22_X1 U1651 ( .A1(n761), .A2(n1774), .B1(n1673), .B2(n1826), .ZN(n2854)
         );
  OAI22_X1 U1652 ( .A1(n762), .A2(n1774), .B1(n1773), .B2(n1827), .ZN(n2853)
         );
  OAI22_X1 U1653 ( .A1(n763), .A2(n1612), .B1(n1673), .B2(n1828), .ZN(n2852)
         );
  OAI22_X1 U1654 ( .A1(n764), .A2(n1774), .B1(n1673), .B2(n1829), .ZN(n2851)
         );
  OAI22_X1 U1655 ( .A1(n765), .A2(n1774), .B1(n1773), .B2(n1830), .ZN(n2850)
         );
  OAI22_X1 U1656 ( .A1(n766), .A2(n1774), .B1(n1773), .B2(n1831), .ZN(n2849)
         );
  OAI22_X1 U1657 ( .A1(n767), .A2(n1774), .B1(n1773), .B2(n1832), .ZN(n2848)
         );
  OAI22_X1 U1658 ( .A1(n768), .A2(n1612), .B1(n1773), .B2(n1833), .ZN(n2847)
         );
  NAND2_X1 U1659 ( .A1(n1776), .A2(n1800), .ZN(n1775) );
  OAI22_X1 U1660 ( .A1(n769), .A2(n1609), .B1(n1777), .B2(n1802), .ZN(n2846)
         );
  OAI22_X1 U1661 ( .A1(n770), .A2(n1609), .B1(n1777), .B2(n1803), .ZN(n2845)
         );
  OAI22_X1 U1662 ( .A1(n771), .A2(n1609), .B1(n1777), .B2(n1804), .ZN(n2844)
         );
  OAI22_X1 U1663 ( .A1(n772), .A2(n1609), .B1(n1777), .B2(n1805), .ZN(n2843)
         );
  OAI22_X1 U1664 ( .A1(n773), .A2(n1609), .B1(n1777), .B2(n1806), .ZN(n2842)
         );
  OAI22_X1 U1665 ( .A1(n774), .A2(n1609), .B1(n1777), .B2(n1807), .ZN(n2841)
         );
  OAI22_X1 U1666 ( .A1(n775), .A2(n1609), .B1(n1777), .B2(n1808), .ZN(n2840)
         );
  OAI22_X1 U1667 ( .A1(n776), .A2(n1609), .B1(n1777), .B2(n1809), .ZN(n2839)
         );
  OAI22_X1 U1668 ( .A1(n777), .A2(n1609), .B1(n1777), .B2(n1810), .ZN(n2838)
         );
  OAI22_X1 U1669 ( .A1(n778), .A2(n1609), .B1(n1777), .B2(n1811), .ZN(n2837)
         );
  OAI22_X1 U1670 ( .A1(n779), .A2(n1609), .B1(n1777), .B2(n1812), .ZN(n2836)
         );
  OAI22_X1 U1671 ( .A1(n780), .A2(n1609), .B1(n1777), .B2(n1813), .ZN(n2835)
         );
  OAI22_X1 U1672 ( .A1(n781), .A2(n1609), .B1(n1674), .B2(n1814), .ZN(n2834)
         );
  OAI22_X1 U1673 ( .A1(n782), .A2(n1609), .B1(n1674), .B2(n1815), .ZN(n2833)
         );
  OAI22_X1 U1674 ( .A1(n783), .A2(n1609), .B1(n1674), .B2(n1816), .ZN(n2832)
         );
  OAI22_X1 U1675 ( .A1(n784), .A2(n1609), .B1(n1674), .B2(n1817), .ZN(n2831)
         );
  OAI22_X1 U1676 ( .A1(n785), .A2(n1609), .B1(n1674), .B2(n1818), .ZN(n2830)
         );
  OAI22_X1 U1677 ( .A1(n786), .A2(n1609), .B1(n1674), .B2(n1819), .ZN(n2829)
         );
  OAI22_X1 U1678 ( .A1(n787), .A2(n1609), .B1(n1674), .B2(n1820), .ZN(n2828)
         );
  OAI22_X1 U1679 ( .A1(n788), .A2(n1609), .B1(n1674), .B2(n1821), .ZN(n2827)
         );
  OAI22_X1 U1680 ( .A1(n789), .A2(n1609), .B1(n1674), .B2(n1822), .ZN(n2826)
         );
  OAI22_X1 U1681 ( .A1(n790), .A2(n1609), .B1(n1674), .B2(n1823), .ZN(n2825)
         );
  OAI22_X1 U1682 ( .A1(n791), .A2(n1609), .B1(n1674), .B2(n1824), .ZN(n2824)
         );
  OAI22_X1 U1683 ( .A1(n792), .A2(n1609), .B1(n1674), .B2(n1825), .ZN(n2823)
         );
  OAI22_X1 U1684 ( .A1(n793), .A2(n1778), .B1(n1777), .B2(n1826), .ZN(n2822)
         );
  OAI22_X1 U1685 ( .A1(n794), .A2(n1778), .B1(n1777), .B2(n1827), .ZN(n2821)
         );
  OAI22_X1 U1686 ( .A1(n795), .A2(n1778), .B1(n1777), .B2(n1828), .ZN(n2820)
         );
  OAI22_X1 U1687 ( .A1(n796), .A2(n1609), .B1(n1674), .B2(n1829), .ZN(n2819)
         );
  OAI22_X1 U1688 ( .A1(n797), .A2(n1778), .B1(n1674), .B2(n1830), .ZN(n2818)
         );
  OAI22_X1 U1689 ( .A1(n798), .A2(n1778), .B1(n1674), .B2(n1831), .ZN(n2817)
         );
  OAI22_X1 U1690 ( .A1(n799), .A2(n1778), .B1(n1674), .B2(n1832), .ZN(n2816)
         );
  OAI22_X1 U1691 ( .A1(n800), .A2(n1609), .B1(n1674), .B2(n1833), .ZN(n2815)
         );
  NAND2_X1 U1692 ( .A1(n1780), .A2(n1800), .ZN(n1779) );
  NAND3_X1 U1693 ( .A1(rst), .A2(n1780), .A3(n1800), .ZN(n1781) );
  OAI22_X1 U1694 ( .A1(n801), .A2(n1584), .B1(n1617), .B2(n1802), .ZN(n2814)
         );
  OAI22_X1 U1695 ( .A1(n802), .A2(n1584), .B1(n1617), .B2(n1803), .ZN(n2813)
         );
  OAI22_X1 U1696 ( .A1(n803), .A2(n1584), .B1(n1617), .B2(n1804), .ZN(n2812)
         );
  OAI22_X1 U1697 ( .A1(n804), .A2(n1584), .B1(n1617), .B2(n1805), .ZN(n2811)
         );
  OAI22_X1 U1698 ( .A1(n805), .A2(n1584), .B1(n1617), .B2(n1806), .ZN(n2810)
         );
  OAI22_X1 U1699 ( .A1(n806), .A2(n1584), .B1(n1617), .B2(n1807), .ZN(n2809)
         );
  OAI22_X1 U1700 ( .A1(n807), .A2(n1584), .B1(n1617), .B2(n1808), .ZN(n2808)
         );
  OAI22_X1 U1701 ( .A1(n808), .A2(n1584), .B1(n1617), .B2(n1809), .ZN(n2807)
         );
  OAI22_X1 U1702 ( .A1(n809), .A2(n1584), .B1(n1617), .B2(n1810), .ZN(n2806)
         );
  OAI22_X1 U1703 ( .A1(n810), .A2(n1584), .B1(n1617), .B2(n1811), .ZN(n2805)
         );
  OAI22_X1 U1704 ( .A1(n811), .A2(n1584), .B1(n1617), .B2(n1812), .ZN(n2804)
         );
  OAI22_X1 U1705 ( .A1(n812), .A2(n1584), .B1(n1617), .B2(n1813), .ZN(n2803)
         );
  OAI22_X1 U1706 ( .A1(n813), .A2(n1584), .B1(n1617), .B2(n1814), .ZN(n2802)
         );
  OAI22_X1 U1707 ( .A1(n814), .A2(n1584), .B1(n1617), .B2(n1815), .ZN(n2801)
         );
  OAI22_X1 U1708 ( .A1(n815), .A2(n1584), .B1(n1617), .B2(n1816), .ZN(n2800)
         );
  OAI22_X1 U1709 ( .A1(n816), .A2(n1584), .B1(n1617), .B2(n1817), .ZN(n2799)
         );
  OAI22_X1 U1710 ( .A1(n817), .A2(n1584), .B1(n1617), .B2(n1818), .ZN(n2798)
         );
  OAI22_X1 U1711 ( .A1(n818), .A2(n1584), .B1(n1617), .B2(n1819), .ZN(n2797)
         );
  OAI22_X1 U1712 ( .A1(n819), .A2(n1584), .B1(n1617), .B2(n1820), .ZN(n2796)
         );
  OAI22_X1 U1713 ( .A1(n820), .A2(n1584), .B1(n1617), .B2(n1821), .ZN(n2795)
         );
  OAI22_X1 U1714 ( .A1(n821), .A2(n1584), .B1(n1617), .B2(n1822), .ZN(n2794)
         );
  OAI22_X1 U1715 ( .A1(n822), .A2(n1584), .B1(n1617), .B2(n1823), .ZN(n2793)
         );
  OAI22_X1 U1716 ( .A1(n823), .A2(n1584), .B1(n1617), .B2(n1824), .ZN(n2792)
         );
  OAI22_X1 U1717 ( .A1(n824), .A2(n1584), .B1(n1617), .B2(n1825), .ZN(n2791)
         );
  OAI22_X1 U1718 ( .A1(n825), .A2(n1782), .B1(n1781), .B2(n1826), .ZN(n2790)
         );
  OAI22_X1 U1719 ( .A1(n826), .A2(n1782), .B1(n1781), .B2(n1827), .ZN(n2789)
         );
  OAI22_X1 U1720 ( .A1(n827), .A2(n1782), .B1(n1781), .B2(n1828), .ZN(n2788)
         );
  OAI22_X1 U1721 ( .A1(n828), .A2(n1584), .B1(n1617), .B2(n1829), .ZN(n2787)
         );
  OAI22_X1 U1722 ( .A1(n829), .A2(n1782), .B1(n1781), .B2(n1830), .ZN(n2786)
         );
  OAI22_X1 U1723 ( .A1(n830), .A2(n1782), .B1(n1617), .B2(n1831), .ZN(n2785)
         );
  OAI22_X1 U1724 ( .A1(n831), .A2(n1782), .B1(n1617), .B2(n1832), .ZN(n2784)
         );
  OAI22_X1 U1725 ( .A1(n832), .A2(n1584), .B1(n1617), .B2(n1833), .ZN(n2783)
         );
  NAND2_X1 U1726 ( .A1(n1784), .A2(n1800), .ZN(n1783) );
  NAND3_X1 U1727 ( .A1(rst), .A2(n1784), .A3(n1800), .ZN(n1785) );
  OAI22_X1 U1728 ( .A1(n833), .A2(n1606), .B1(n1621), .B2(n1802), .ZN(n2782)
         );
  OAI22_X1 U1729 ( .A1(n834), .A2(n1606), .B1(n1621), .B2(n1803), .ZN(n2781)
         );
  OAI22_X1 U1730 ( .A1(n835), .A2(n1606), .B1(n1621), .B2(n1804), .ZN(n2780)
         );
  OAI22_X1 U1731 ( .A1(n836), .A2(n1606), .B1(n1621), .B2(n1805), .ZN(n2779)
         );
  OAI22_X1 U1732 ( .A1(n837), .A2(n1606), .B1(n1621), .B2(n1806), .ZN(n2778)
         );
  OAI22_X1 U1733 ( .A1(n838), .A2(n1606), .B1(n1621), .B2(n1807), .ZN(n2777)
         );
  OAI22_X1 U1734 ( .A1(n839), .A2(n1606), .B1(n1621), .B2(n1808), .ZN(n2776)
         );
  OAI22_X1 U1735 ( .A1(n840), .A2(n1606), .B1(n1621), .B2(n1809), .ZN(n2775)
         );
  OAI22_X1 U1736 ( .A1(n841), .A2(n1606), .B1(n1621), .B2(n1810), .ZN(n2774)
         );
  OAI22_X1 U1737 ( .A1(n842), .A2(n1606), .B1(n1621), .B2(n1811), .ZN(n2773)
         );
  OAI22_X1 U1738 ( .A1(n843), .A2(n1606), .B1(n1621), .B2(n1812), .ZN(n2772)
         );
  OAI22_X1 U1739 ( .A1(n844), .A2(n1606), .B1(n1621), .B2(n1813), .ZN(n2771)
         );
  OAI22_X1 U1740 ( .A1(n845), .A2(n1606), .B1(n1621), .B2(n1814), .ZN(n2770)
         );
  OAI22_X1 U1741 ( .A1(n846), .A2(n1606), .B1(n1621), .B2(n1815), .ZN(n2769)
         );
  OAI22_X1 U1742 ( .A1(n847), .A2(n1606), .B1(n1621), .B2(n1816), .ZN(n2768)
         );
  OAI22_X1 U1743 ( .A1(n848), .A2(n1606), .B1(n1621), .B2(n1817), .ZN(n2767)
         );
  OAI22_X1 U1744 ( .A1(n849), .A2(n1606), .B1(n1621), .B2(n1818), .ZN(n2766)
         );
  OAI22_X1 U1745 ( .A1(n850), .A2(n1606), .B1(n1621), .B2(n1819), .ZN(n2765)
         );
  OAI22_X1 U1746 ( .A1(n851), .A2(n1606), .B1(n1621), .B2(n1820), .ZN(n2764)
         );
  OAI22_X1 U1747 ( .A1(n852), .A2(n1606), .B1(n1621), .B2(n1821), .ZN(n2763)
         );
  OAI22_X1 U1748 ( .A1(n853), .A2(n1606), .B1(n1621), .B2(n1822), .ZN(n2762)
         );
  OAI22_X1 U1749 ( .A1(n854), .A2(n1606), .B1(n1621), .B2(n1823), .ZN(n2761)
         );
  OAI22_X1 U1750 ( .A1(n855), .A2(n1606), .B1(n1621), .B2(n1824), .ZN(n2760)
         );
  OAI22_X1 U1751 ( .A1(n856), .A2(n1606), .B1(n1621), .B2(n1825), .ZN(n2759)
         );
  OAI22_X1 U1752 ( .A1(n857), .A2(n1786), .B1(n1785), .B2(n1826), .ZN(n2758)
         );
  OAI22_X1 U1753 ( .A1(n858), .A2(n1786), .B1(n1785), .B2(n1827), .ZN(n2757)
         );
  OAI22_X1 U1754 ( .A1(n859), .A2(n1786), .B1(n1785), .B2(n1828), .ZN(n2756)
         );
  OAI22_X1 U1755 ( .A1(n860), .A2(n1606), .B1(n1621), .B2(n1829), .ZN(n2755)
         );
  OAI22_X1 U1756 ( .A1(n861), .A2(n1786), .B1(n1785), .B2(n1830), .ZN(n2754)
         );
  OAI22_X1 U1757 ( .A1(n862), .A2(n1786), .B1(n1621), .B2(n1831), .ZN(n2753)
         );
  OAI22_X1 U1758 ( .A1(n863), .A2(n1786), .B1(n1621), .B2(n1832), .ZN(n2752)
         );
  OAI22_X1 U1759 ( .A1(n864), .A2(n1606), .B1(n1621), .B2(n1833), .ZN(n2751)
         );
  NAND2_X1 U1760 ( .A1(n1788), .A2(n1800), .ZN(n1787) );
  OAI22_X1 U1761 ( .A1(n865), .A2(n1601), .B1(n1789), .B2(n1802), .ZN(n2750)
         );
  OAI22_X1 U1762 ( .A1(n866), .A2(n1601), .B1(n1789), .B2(n1803), .ZN(n2749)
         );
  OAI22_X1 U1763 ( .A1(n867), .A2(n1601), .B1(n1789), .B2(n1804), .ZN(n2748)
         );
  OAI22_X1 U1764 ( .A1(n868), .A2(n1601), .B1(n1789), .B2(n1805), .ZN(n2747)
         );
  OAI22_X1 U1765 ( .A1(n869), .A2(n1601), .B1(n1789), .B2(n1806), .ZN(n2746)
         );
  OAI22_X1 U1766 ( .A1(n870), .A2(n1601), .B1(n1789), .B2(n1807), .ZN(n2745)
         );
  OAI22_X1 U1767 ( .A1(n871), .A2(n1601), .B1(n1789), .B2(n1808), .ZN(n2744)
         );
  OAI22_X1 U1768 ( .A1(n872), .A2(n1601), .B1(n1789), .B2(n1809), .ZN(n2743)
         );
  OAI22_X1 U1769 ( .A1(n873), .A2(n1601), .B1(n1789), .B2(n1810), .ZN(n2742)
         );
  OAI22_X1 U1770 ( .A1(n874), .A2(n1601), .B1(n1789), .B2(n1811), .ZN(n2741)
         );
  OAI22_X1 U1771 ( .A1(n875), .A2(n1601), .B1(n1789), .B2(n1812), .ZN(n2740)
         );
  OAI22_X1 U1772 ( .A1(n876), .A2(n1601), .B1(n1789), .B2(n1813), .ZN(n2739)
         );
  OAI22_X1 U1773 ( .A1(n877), .A2(n1601), .B1(n1675), .B2(n1814), .ZN(n2738)
         );
  OAI22_X1 U1774 ( .A1(n878), .A2(n1601), .B1(n1675), .B2(n1815), .ZN(n2737)
         );
  OAI22_X1 U1775 ( .A1(n879), .A2(n1601), .B1(n1675), .B2(n1816), .ZN(n2736)
         );
  OAI22_X1 U1776 ( .A1(n880), .A2(n1601), .B1(n1675), .B2(n1817), .ZN(n2735)
         );
  OAI22_X1 U1777 ( .A1(n881), .A2(n1601), .B1(n1675), .B2(n1818), .ZN(n2734)
         );
  OAI22_X1 U1778 ( .A1(n882), .A2(n1601), .B1(n1675), .B2(n1819), .ZN(n2733)
         );
  OAI22_X1 U1779 ( .A1(n883), .A2(n1601), .B1(n1675), .B2(n1820), .ZN(n2732)
         );
  OAI22_X1 U1780 ( .A1(n884), .A2(n1601), .B1(n1675), .B2(n1821), .ZN(n2731)
         );
  OAI22_X1 U1781 ( .A1(n885), .A2(n1601), .B1(n1675), .B2(n1822), .ZN(n2730)
         );
  OAI22_X1 U1782 ( .A1(n886), .A2(n1601), .B1(n1675), .B2(n1823), .ZN(n2729)
         );
  OAI22_X1 U1783 ( .A1(n887), .A2(n1601), .B1(n1675), .B2(n1824), .ZN(n2728)
         );
  OAI22_X1 U1784 ( .A1(n888), .A2(n1601), .B1(n1675), .B2(n1825), .ZN(n2727)
         );
  OAI22_X1 U1785 ( .A1(n889), .A2(n1790), .B1(n1789), .B2(n1826), .ZN(n2726)
         );
  OAI22_X1 U1786 ( .A1(n890), .A2(n1790), .B1(n1789), .B2(n1827), .ZN(n2725)
         );
  OAI22_X1 U1787 ( .A1(n891), .A2(n1790), .B1(n1789), .B2(n1828), .ZN(n2724)
         );
  OAI22_X1 U1788 ( .A1(n892), .A2(n1601), .B1(n1675), .B2(n1829), .ZN(n2723)
         );
  OAI22_X1 U1789 ( .A1(n893), .A2(n1790), .B1(n1675), .B2(n1830), .ZN(n2722)
         );
  OAI22_X1 U1790 ( .A1(n894), .A2(n1790), .B1(n1675), .B2(n1831), .ZN(n2721)
         );
  OAI22_X1 U1791 ( .A1(n895), .A2(n1790), .B1(n1675), .B2(n1832), .ZN(n2720)
         );
  OAI22_X1 U1792 ( .A1(n896), .A2(n1601), .B1(n1675), .B2(n1833), .ZN(n2719)
         );
  NAND2_X1 U1793 ( .A1(n1792), .A2(n1800), .ZN(n1791) );
  OAI22_X1 U1794 ( .A1(n897), .A2(n1596), .B1(n1793), .B2(n1802), .ZN(n2718)
         );
  OAI22_X1 U1795 ( .A1(n898), .A2(n1596), .B1(n1793), .B2(n1803), .ZN(n2717)
         );
  OAI22_X1 U1796 ( .A1(n899), .A2(n1596), .B1(n1793), .B2(n1804), .ZN(n2716)
         );
  OAI22_X1 U1797 ( .A1(n900), .A2(n1596), .B1(n1793), .B2(n1805), .ZN(n2715)
         );
  OAI22_X1 U1798 ( .A1(n901), .A2(n1596), .B1(n1793), .B2(n1806), .ZN(n2714)
         );
  OAI22_X1 U1799 ( .A1(n902), .A2(n1596), .B1(n1793), .B2(n1807), .ZN(n2713)
         );
  OAI22_X1 U1800 ( .A1(n903), .A2(n1596), .B1(n1793), .B2(n1808), .ZN(n2712)
         );
  OAI22_X1 U1801 ( .A1(n904), .A2(n1596), .B1(n1793), .B2(n1809), .ZN(n2711)
         );
  OAI22_X1 U1802 ( .A1(n905), .A2(n1596), .B1(n1793), .B2(n1810), .ZN(n2710)
         );
  OAI22_X1 U1803 ( .A1(n906), .A2(n1596), .B1(n1793), .B2(n1811), .ZN(n2709)
         );
  OAI22_X1 U1804 ( .A1(n907), .A2(n1596), .B1(n1793), .B2(n1812), .ZN(n2708)
         );
  OAI22_X1 U1805 ( .A1(n908), .A2(n1596), .B1(n1793), .B2(n1813), .ZN(n2707)
         );
  OAI22_X1 U1806 ( .A1(n909), .A2(n1596), .B1(n1676), .B2(n1814), .ZN(n2706)
         );
  OAI22_X1 U1807 ( .A1(n910), .A2(n1596), .B1(n1676), .B2(n1815), .ZN(n2705)
         );
  OAI22_X1 U1808 ( .A1(n911), .A2(n1596), .B1(n1676), .B2(n1816), .ZN(n2704)
         );
  OAI22_X1 U1809 ( .A1(n912), .A2(n1596), .B1(n1676), .B2(n1817), .ZN(n2703)
         );
  OAI22_X1 U1810 ( .A1(n913), .A2(n1596), .B1(n1676), .B2(n1818), .ZN(n2702)
         );
  OAI22_X1 U1811 ( .A1(n914), .A2(n1596), .B1(n1676), .B2(n1819), .ZN(n2701)
         );
  OAI22_X1 U1812 ( .A1(n915), .A2(n1596), .B1(n1676), .B2(n1820), .ZN(n2700)
         );
  OAI22_X1 U1813 ( .A1(n916), .A2(n1596), .B1(n1676), .B2(n1821), .ZN(n2699)
         );
  OAI22_X1 U1814 ( .A1(n917), .A2(n1596), .B1(n1676), .B2(n1822), .ZN(n2698)
         );
  OAI22_X1 U1815 ( .A1(n918), .A2(n1596), .B1(n1676), .B2(n1823), .ZN(n2697)
         );
  OAI22_X1 U1816 ( .A1(n919), .A2(n1596), .B1(n1676), .B2(n1824), .ZN(n2696)
         );
  OAI22_X1 U1817 ( .A1(n920), .A2(n1596), .B1(n1676), .B2(n1825), .ZN(n2695)
         );
  OAI22_X1 U1818 ( .A1(n921), .A2(n1794), .B1(n1793), .B2(n1826), .ZN(n2694)
         );
  OAI22_X1 U1819 ( .A1(n922), .A2(n1794), .B1(n1793), .B2(n1827), .ZN(n2693)
         );
  OAI22_X1 U1820 ( .A1(n923), .A2(n1794), .B1(n1793), .B2(n1828), .ZN(n2692)
         );
  OAI22_X1 U1821 ( .A1(n924), .A2(n1596), .B1(n1676), .B2(n1829), .ZN(n2691)
         );
  OAI22_X1 U1822 ( .A1(n925), .A2(n1794), .B1(n1676), .B2(n1830), .ZN(n2690)
         );
  OAI22_X1 U1823 ( .A1(n926), .A2(n1794), .B1(n1676), .B2(n1831), .ZN(n2689)
         );
  OAI22_X1 U1824 ( .A1(n927), .A2(n1794), .B1(n1676), .B2(n1832), .ZN(n2688)
         );
  OAI22_X1 U1825 ( .A1(n928), .A2(n1596), .B1(n1676), .B2(n1833), .ZN(n2687)
         );
  NAND2_X1 U1826 ( .A1(n1796), .A2(n1800), .ZN(n1795) );
  NAND3_X1 U1827 ( .A1(rst), .A2(n1796), .A3(n1800), .ZN(n1797) );
  OAI22_X1 U1828 ( .A1(n929), .A2(n1586), .B1(n1616), .B2(n1802), .ZN(n2686)
         );
  OAI22_X1 U1829 ( .A1(n930), .A2(n1586), .B1(n1616), .B2(n1803), .ZN(n2685)
         );
  OAI22_X1 U1830 ( .A1(n931), .A2(n1586), .B1(n1616), .B2(n1804), .ZN(n2684)
         );
  OAI22_X1 U1831 ( .A1(n932), .A2(n1586), .B1(n1616), .B2(n1805), .ZN(n2683)
         );
  OAI22_X1 U1832 ( .A1(n933), .A2(n1586), .B1(n1616), .B2(n1806), .ZN(n2682)
         );
  OAI22_X1 U1833 ( .A1(n934), .A2(n1586), .B1(n1616), .B2(n1807), .ZN(n2681)
         );
  OAI22_X1 U1834 ( .A1(n935), .A2(n1586), .B1(n1616), .B2(n1808), .ZN(n2680)
         );
  OAI22_X1 U1835 ( .A1(n936), .A2(n1586), .B1(n1616), .B2(n1809), .ZN(n2679)
         );
  OAI22_X1 U1836 ( .A1(n937), .A2(n1586), .B1(n1616), .B2(n1810), .ZN(n2678)
         );
  OAI22_X1 U1837 ( .A1(n938), .A2(n1586), .B1(n1616), .B2(n1811), .ZN(n2677)
         );
  OAI22_X1 U1838 ( .A1(n939), .A2(n1586), .B1(n1616), .B2(n1812), .ZN(n2676)
         );
  OAI22_X1 U1839 ( .A1(n940), .A2(n1586), .B1(n1616), .B2(n1813), .ZN(n2675)
         );
  OAI22_X1 U1840 ( .A1(n941), .A2(n1586), .B1(n1616), .B2(n1814), .ZN(n2674)
         );
  OAI22_X1 U1841 ( .A1(n942), .A2(n1586), .B1(n1616), .B2(n1815), .ZN(n2673)
         );
  OAI22_X1 U1842 ( .A1(n943), .A2(n1586), .B1(n1616), .B2(n1816), .ZN(n2672)
         );
  OAI22_X1 U1843 ( .A1(n944), .A2(n1586), .B1(n1616), .B2(n1817), .ZN(n2671)
         );
  OAI22_X1 U1844 ( .A1(n945), .A2(n1586), .B1(n1616), .B2(n1818), .ZN(n2670)
         );
  OAI22_X1 U1845 ( .A1(n946), .A2(n1586), .B1(n1616), .B2(n1819), .ZN(n2669)
         );
  OAI22_X1 U1846 ( .A1(n947), .A2(n1586), .B1(n1616), .B2(n1820), .ZN(n2668)
         );
  OAI22_X1 U1847 ( .A1(n948), .A2(n1586), .B1(n1616), .B2(n1821), .ZN(n2667)
         );
  OAI22_X1 U1848 ( .A1(n949), .A2(n1586), .B1(n1616), .B2(n1822), .ZN(n2666)
         );
  OAI22_X1 U1849 ( .A1(n950), .A2(n1586), .B1(n1616), .B2(n1823), .ZN(n2665)
         );
  OAI22_X1 U1850 ( .A1(n951), .A2(n1586), .B1(n1616), .B2(n1824), .ZN(n2664)
         );
  OAI22_X1 U1851 ( .A1(n952), .A2(n1586), .B1(n1616), .B2(n1825), .ZN(n2663)
         );
  OAI22_X1 U1852 ( .A1(n953), .A2(n1798), .B1(n1616), .B2(n1826), .ZN(n2662)
         );
  OAI22_X1 U1853 ( .A1(n954), .A2(n1586), .B1(n1616), .B2(n1827), .ZN(n2661)
         );
  OAI22_X1 U1854 ( .A1(n955), .A2(n1798), .B1(n1616), .B2(n1828), .ZN(n2660)
         );
  OAI22_X1 U1855 ( .A1(n956), .A2(n1586), .B1(n1616), .B2(n1829), .ZN(n2659)
         );
  OAI22_X1 U1856 ( .A1(n957), .A2(n1798), .B1(n1797), .B2(n1830), .ZN(n2658)
         );
  OAI22_X1 U1857 ( .A1(n958), .A2(n1798), .B1(n1797), .B2(n1831), .ZN(n2657)
         );
  OAI22_X1 U1858 ( .A1(n959), .A2(n1798), .B1(n1797), .B2(n1832), .ZN(n2656)
         );
  OAI22_X1 U1859 ( .A1(n960), .A2(n1798), .B1(n1797), .B2(n1833), .ZN(n2655)
         );
  NAND2_X1 U1860 ( .A1(n1801), .A2(n1800), .ZN(n1799) );
  NAND3_X1 U1861 ( .A1(rst), .A2(n1801), .A3(n1800), .ZN(n1834) );
  OAI22_X1 U1862 ( .A1(n961), .A2(n1592), .B1(n1620), .B2(n1802), .ZN(n2654)
         );
  OAI22_X1 U1863 ( .A1(n962), .A2(n1592), .B1(n1620), .B2(n1803), .ZN(n2653)
         );
  OAI22_X1 U1864 ( .A1(n963), .A2(n1592), .B1(n1620), .B2(n1804), .ZN(n2652)
         );
  OAI22_X1 U1865 ( .A1(n964), .A2(n1592), .B1(n1620), .B2(n1805), .ZN(n2651)
         );
  OAI22_X1 U1866 ( .A1(n965), .A2(n1592), .B1(n1620), .B2(n1806), .ZN(n2650)
         );
  OAI22_X1 U1867 ( .A1(n966), .A2(n1592), .B1(n1620), .B2(n1807), .ZN(n2649)
         );
  OAI22_X1 U1868 ( .A1(n967), .A2(n1592), .B1(n1620), .B2(n1808), .ZN(n2648)
         );
  OAI22_X1 U1869 ( .A1(n968), .A2(n1592), .B1(n1620), .B2(n1809), .ZN(n2647)
         );
  OAI22_X1 U1870 ( .A1(n969), .A2(n1592), .B1(n1620), .B2(n1810), .ZN(n2646)
         );
  OAI22_X1 U1871 ( .A1(n970), .A2(n1592), .B1(n1620), .B2(n1811), .ZN(n2645)
         );
  OAI22_X1 U1872 ( .A1(n971), .A2(n1592), .B1(n1620), .B2(n1812), .ZN(n2644)
         );
  OAI22_X1 U1873 ( .A1(n972), .A2(n1592), .B1(n1620), .B2(n1813), .ZN(n2643)
         );
  OAI22_X1 U1874 ( .A1(n973), .A2(n1592), .B1(n1620), .B2(n1814), .ZN(n2642)
         );
  OAI22_X1 U1875 ( .A1(n974), .A2(n1592), .B1(n1620), .B2(n1815), .ZN(n2641)
         );
  OAI22_X1 U1876 ( .A1(n975), .A2(n1592), .B1(n1620), .B2(n1816), .ZN(n2640)
         );
  OAI22_X1 U1877 ( .A1(n976), .A2(n1592), .B1(n1620), .B2(n1817), .ZN(n2639)
         );
  OAI22_X1 U1878 ( .A1(n977), .A2(n1592), .B1(n1620), .B2(n1818), .ZN(n2638)
         );
  OAI22_X1 U1879 ( .A1(n978), .A2(n1592), .B1(n1620), .B2(n1819), .ZN(n2637)
         );
  OAI22_X1 U1880 ( .A1(n979), .A2(n1592), .B1(n1620), .B2(n1820), .ZN(n2636)
         );
  OAI22_X1 U1881 ( .A1(n980), .A2(n1592), .B1(n1620), .B2(n1821), .ZN(n2635)
         );
  OAI22_X1 U1882 ( .A1(n981), .A2(n1592), .B1(n1620), .B2(n1822), .ZN(n2634)
         );
  OAI22_X1 U1883 ( .A1(n982), .A2(n1592), .B1(n1620), .B2(n1823), .ZN(n2633)
         );
  OAI22_X1 U1884 ( .A1(n983), .A2(n1592), .B1(n1620), .B2(n1824), .ZN(n2632)
         );
  OAI22_X1 U1885 ( .A1(n984), .A2(n1592), .B1(n1620), .B2(n1825), .ZN(n2631)
         );
  OAI22_X1 U1886 ( .A1(n985), .A2(n1835), .B1(n1620), .B2(n1826), .ZN(n2630)
         );
  OAI22_X1 U1887 ( .A1(n986), .A2(n1592), .B1(n1620), .B2(n1827), .ZN(n2629)
         );
  OAI22_X1 U1888 ( .A1(n987), .A2(n1592), .B1(n1620), .B2(n1828), .ZN(n2628)
         );
  OAI22_X1 U1889 ( .A1(n988), .A2(n1835), .B1(n1620), .B2(n1829), .ZN(n2627)
         );
  OAI22_X1 U1890 ( .A1(n989), .A2(n1835), .B1(n1834), .B2(n1830), .ZN(n2626)
         );
  OAI22_X1 U1891 ( .A1(n990), .A2(n1835), .B1(n1834), .B2(n1831), .ZN(n2625)
         );
  OAI22_X1 U1892 ( .A1(n991), .A2(n1835), .B1(n1834), .B2(n1832), .ZN(n2624)
         );
  OAI22_X1 U1893 ( .A1(n992), .A2(n1835), .B1(n1834), .B2(n1833), .ZN(n2623)
         );
  OAI221_X1 U1894 ( .B1(n1686), .B2(lo_out[0]), .C1(n1688), .C2(lo_in[0]), .A(
        rst), .ZN(n2547) );
  OAI221_X1 U1895 ( .B1(n1686), .B2(lo_out[1]), .C1(n1688), .C2(lo_in[1]), .A(
        rst), .ZN(n2546) );
  OAI221_X1 U1896 ( .B1(n1686), .B2(lo_out[2]), .C1(n1688), .C2(lo_in[2]), .A(
        rst), .ZN(n2545) );
  OAI221_X1 U1897 ( .B1(n1686), .B2(lo_out[3]), .C1(n1688), .C2(lo_in[3]), .A(
        rst), .ZN(n2544) );
  OAI221_X1 U1898 ( .B1(n1686), .B2(lo_out[4]), .C1(n1688), .C2(lo_in[4]), .A(
        rst), .ZN(n2543) );
  OAI221_X1 U1899 ( .B1(n1686), .B2(lo_out[5]), .C1(n1688), .C2(lo_in[5]), .A(
        rst), .ZN(n2542) );
  OAI221_X1 U1900 ( .B1(n1686), .B2(lo_out[6]), .C1(n1688), .C2(lo_in[6]), .A(
        rst), .ZN(n2541) );
  OAI221_X1 U1901 ( .B1(n1686), .B2(lo_out[7]), .C1(n1688), .C2(lo_in[7]), .A(
        rst), .ZN(n2540) );
  OAI221_X1 U1902 ( .B1(n1686), .B2(lo_out[8]), .C1(n1615), .C2(lo_in[8]), .A(
        rst), .ZN(n2539) );
  OAI221_X1 U1903 ( .B1(n1686), .B2(lo_out[9]), .C1(n1615), .C2(lo_in[9]), .A(
        rst), .ZN(n2538) );
  OAI221_X1 U1904 ( .B1(n1686), .B2(lo_out[10]), .C1(n1615), .C2(lo_in[10]), 
        .A(rst), .ZN(n2537) );
  OAI221_X1 U1905 ( .B1(n1686), .B2(lo_out[11]), .C1(n1615), .C2(lo_in[11]), 
        .A(rst), .ZN(n2536) );
  OAI221_X1 U1906 ( .B1(hilo_wr_en), .B2(lo_out[12]), .C1(n1615), .C2(
        lo_in[12]), .A(rst), .ZN(n2535) );
  OAI221_X1 U1907 ( .B1(hilo_wr_en), .B2(lo_out[13]), .C1(n1615), .C2(
        lo_in[13]), .A(rst), .ZN(n2534) );
  OAI221_X1 U1908 ( .B1(hilo_wr_en), .B2(lo_out[14]), .C1(n1615), .C2(
        lo_in[14]), .A(rst), .ZN(n2533) );
  OAI221_X1 U1909 ( .B1(hilo_wr_en), .B2(lo_out[15]), .C1(n1622), .C2(
        lo_in[15]), .A(rst), .ZN(n2532) );
  OAI221_X1 U1910 ( .B1(hilo_wr_en), .B2(lo_out[16]), .C1(n1622), .C2(
        lo_in[16]), .A(rst), .ZN(n2531) );
  OAI221_X1 U1911 ( .B1(hilo_wr_en), .B2(lo_out[17]), .C1(n1622), .C2(
        lo_in[17]), .A(rst), .ZN(n2530) );
  OAI221_X1 U1912 ( .B1(n1686), .B2(lo_out[18]), .C1(n1622), .C2(lo_in[18]), 
        .A(rst), .ZN(n2529) );
  OAI221_X1 U1913 ( .B1(n1687), .B2(lo_out[19]), .C1(n1622), .C2(lo_in[19]), 
        .A(rst), .ZN(n2528) );
  OAI221_X1 U1914 ( .B1(n1687), .B2(lo_out[20]), .C1(n1622), .C2(lo_in[20]), 
        .A(rst), .ZN(n2527) );
  OAI221_X1 U1915 ( .B1(n1686), .B2(lo_out[21]), .C1(n1622), .C2(lo_in[21]), 
        .A(rst), .ZN(n2526) );
  OAI221_X1 U1916 ( .B1(hilo_wr_en), .B2(lo_out[22]), .C1(n1688), .C2(
        lo_in[22]), .A(rst), .ZN(n2525) );
  OAI221_X1 U1917 ( .B1(n1687), .B2(lo_out[23]), .C1(n1615), .C2(lo_in[23]), 
        .A(rst), .ZN(n2524) );
  OAI221_X1 U1918 ( .B1(n1687), .B2(lo_out[24]), .C1(n1688), .C2(lo_in[24]), 
        .A(rst), .ZN(n2523) );
  OAI221_X1 U1919 ( .B1(n1687), .B2(lo_out[25]), .C1(n1622), .C2(lo_in[25]), 
        .A(rst), .ZN(n2522) );
  OAI221_X1 U1920 ( .B1(n1687), .B2(lo_out[26]), .C1(n1688), .C2(lo_in[26]), 
        .A(rst), .ZN(n2521) );
  OAI221_X1 U1921 ( .B1(n1687), .B2(lo_out[27]), .C1(n1582), .C2(lo_in[27]), 
        .A(rst), .ZN(n2520) );
  OAI221_X1 U1922 ( .B1(n1687), .B2(lo_out[28]), .C1(n1688), .C2(lo_in[28]), 
        .A(rst), .ZN(n2519) );
  OAI221_X1 U1923 ( .B1(n1687), .B2(lo_out[29]), .C1(n1615), .C2(lo_in[29]), 
        .A(rst), .ZN(n2518) );
  OAI221_X1 U1924 ( .B1(n1687), .B2(lo_out[30]), .C1(n1615), .C2(lo_in[30]), 
        .A(rst), .ZN(n2517) );
  OAI221_X1 U1925 ( .B1(n1687), .B2(lo_out[31]), .C1(n1615), .C2(lo_in[31]), 
        .A(rst), .ZN(n2516) );
  OAI221_X1 U1926 ( .B1(n1687), .B2(hi_out[0]), .C1(n1615), .C2(hi_in[0]), .A(
        rst), .ZN(n2515) );
  OAI221_X1 U1927 ( .B1(n1687), .B2(hi_out[1]), .C1(n1615), .C2(hi_in[1]), .A(
        rst), .ZN(n2514) );
  OAI221_X1 U1928 ( .B1(n1687), .B2(hi_out[2]), .C1(n1615), .C2(hi_in[2]), .A(
        rst), .ZN(n2513) );
  OAI221_X1 U1929 ( .B1(n1687), .B2(hi_out[3]), .C1(n1615), .C2(hi_in[3]), .A(
        rst), .ZN(n2512) );
  OAI221_X1 U1930 ( .B1(n1686), .B2(hi_out[4]), .C1(n1582), .C2(hi_in[4]), .A(
        rst), .ZN(n2511) );
  OAI221_X1 U1931 ( .B1(n1687), .B2(hi_out[5]), .C1(n1582), .C2(hi_in[5]), .A(
        rst), .ZN(n2510) );
  OAI221_X1 U1932 ( .B1(hilo_wr_en), .B2(hi_out[6]), .C1(n1582), .C2(hi_in[6]), 
        .A(rst), .ZN(n2509) );
  OAI221_X1 U1933 ( .B1(n1687), .B2(hi_out[7]), .C1(n1582), .C2(hi_in[7]), .A(
        rst), .ZN(n2508) );
  OAI221_X1 U1934 ( .B1(n1687), .B2(hi_out[8]), .C1(n1582), .C2(hi_in[8]), .A(
        rst), .ZN(n2507) );
  OAI221_X1 U1935 ( .B1(n1686), .B2(hi_out[9]), .C1(n1582), .C2(hi_in[9]), .A(
        rst), .ZN(n2506) );
  OAI221_X1 U1936 ( .B1(n1686), .B2(hi_out[10]), .C1(n1582), .C2(hi_in[10]), 
        .A(rst), .ZN(n2505) );
  OAI221_X1 U1937 ( .B1(hilo_wr_en), .B2(hi_out[11]), .C1(n1688), .C2(
        hi_in[11]), .A(rst), .ZN(n2504) );
  OAI221_X1 U1938 ( .B1(n1686), .B2(hi_out[12]), .C1(n1688), .C2(hi_in[12]), 
        .A(rst), .ZN(n2503) );
  OAI221_X1 U1939 ( .B1(n1687), .B2(hi_out[13]), .C1(n1688), .C2(hi_in[13]), 
        .A(rst), .ZN(n2502) );
  OAI221_X1 U1940 ( .B1(n1687), .B2(hi_out[14]), .C1(n1688), .C2(hi_in[14]), 
        .A(rst), .ZN(n2501) );
  OAI221_X1 U1941 ( .B1(hilo_wr_en), .B2(hi_out[15]), .C1(n1688), .C2(
        hi_in[15]), .A(rst), .ZN(n2500) );
  OAI221_X1 U1942 ( .B1(hilo_wr_en), .B2(hi_out[16]), .C1(n1688), .C2(
        hi_in[16]), .A(rst), .ZN(n2499) );
  OAI221_X1 U1943 ( .B1(hilo_wr_en), .B2(hi_out[17]), .C1(n1688), .C2(
        hi_in[17]), .A(rst), .ZN(n2498) );
  OAI221_X1 U1944 ( .B1(n1686), .B2(hi_out[18]), .C1(n1582), .C2(hi_in[18]), 
        .A(rst), .ZN(n2497) );
  OAI221_X1 U1945 ( .B1(hilo_wr_en), .B2(hi_out[19]), .C1(n1582), .C2(
        hi_in[19]), .A(rst), .ZN(n2496) );
  OAI221_X1 U1946 ( .B1(hilo_wr_en), .B2(hi_out[20]), .C1(n1582), .C2(
        hi_in[20]), .A(rst), .ZN(n2495) );
  OAI221_X1 U1947 ( .B1(hilo_wr_en), .B2(hi_out[21]), .C1(n1582), .C2(
        hi_in[21]), .A(rst), .ZN(n2494) );
  OAI221_X1 U1948 ( .B1(hilo_wr_en), .B2(hi_out[22]), .C1(n1582), .C2(
        hi_in[22]), .A(rst), .ZN(n2493) );
  OAI221_X1 U1949 ( .B1(hilo_wr_en), .B2(hi_out[23]), .C1(n1582), .C2(
        hi_in[23]), .A(rst), .ZN(n2492) );
  OAI221_X1 U1950 ( .B1(hilo_wr_en), .B2(hi_out[24]), .C1(n1582), .C2(
        hi_in[24]), .A(rst), .ZN(n2491) );
  OAI221_X1 U1951 ( .B1(hilo_wr_en), .B2(hi_out[25]), .C1(n1622), .C2(
        hi_in[25]), .A(rst), .ZN(n2490) );
  OAI221_X1 U1952 ( .B1(hilo_wr_en), .B2(hi_out[26]), .C1(n1622), .C2(
        hi_in[26]), .A(rst), .ZN(n2489) );
  OAI221_X1 U1953 ( .B1(hilo_wr_en), .B2(hi_out[27]), .C1(n1622), .C2(
        hi_in[27]), .A(rst), .ZN(n2488) );
  OAI221_X1 U1954 ( .B1(hilo_wr_en), .B2(hi_out[28]), .C1(n1622), .C2(
        hi_in[28]), .A(rst), .ZN(n2487) );
  OAI221_X1 U1955 ( .B1(n1686), .B2(hi_out[29]), .C1(n1622), .C2(hi_in[29]), 
        .A(rst), .ZN(n2486) );
  OAI221_X1 U1956 ( .B1(n1687), .B2(hi_out[30]), .C1(n1622), .C2(hi_in[30]), 
        .A(rst), .ZN(n2485) );
  OAI221_X1 U1957 ( .B1(n1686), .B2(hi_out[31]), .C1(n1622), .C2(hi_in[31]), 
        .A(rst), .ZN(n2482) );
  INV_X1 U1958 ( .A(rp1_out_sel[0]), .ZN(n1853) );
  NOR2_X1 U1959 ( .A1(rp1_out_sel[1]), .A2(rp1_out_sel[0]), .ZN(n2282) );
  INV_X1 U1960 ( .A(rp1_addr[2]), .ZN(n1836) );
  NOR2_X1 U1961 ( .A1(rp1_addr[1]), .A2(n1836), .ZN(n1847) );
  INV_X1 U1962 ( .A(rp1_addr[4]), .ZN(n1841) );
  NOR3_X1 U1963 ( .A1(rp1_addr[0]), .A2(rp1_addr[3]), .A3(n1841), .ZN(n1842)
         );
  NAND2_X1 U1964 ( .A1(n1847), .A2(n1842), .ZN(n2271) );
  NAND2_X1 U1965 ( .A1(rp1_addr[4]), .A2(rp1_addr[3]), .ZN(n1837) );
  NOR2_X1 U1966 ( .A1(rp1_addr[0]), .A2(n1837), .ZN(n1839) );
  NOR2_X1 U1967 ( .A1(rp1_addr[2]), .A2(rp1_addr[1]), .ZN(n1845) );
  AND2_X1 U1968 ( .A1(rp1_addr[2]), .A2(rp1_addr[1]), .ZN(n1852) );
  INV_X1 U1969 ( .A(rp1_addr[0]), .ZN(n1840) );
  INV_X1 U1970 ( .A(rp1_addr[3]), .ZN(n1838) );
  NOR3_X1 U1971 ( .A1(rp1_addr[4]), .A2(n1840), .A3(n1838), .ZN(n1843) );
  AND2_X1 U1972 ( .A1(n1836), .A2(rp1_addr[1]), .ZN(n1850) );
  NOR2_X1 U1973 ( .A1(n1840), .A2(n1837), .ZN(n1844) );
  NOR3_X1 U1974 ( .A1(rp1_addr[0]), .A2(rp1_addr[4]), .A3(n1838), .ZN(n1851)
         );
  NOR3_X1 U1975 ( .A1(rp1_addr[4]), .A2(rp1_addr[3]), .A3(n1840), .ZN(n1846)
         );
  NOR3_X1 U1976 ( .A1(rp1_addr[3]), .A2(n1841), .A3(n1840), .ZN(n1848) );
  NOR3_X1 U1977 ( .A1(rp1_addr[0]), .A2(rp1_addr[4]), .A3(rp1_addr[3]), .ZN(
        n1849) );
  NAND2_X1 U1978 ( .A1(n1847), .A2(n1846), .ZN(n2254) );
  NOR2_X1 U1979 ( .A1(rp1_out_sel[1]), .A2(n1853), .ZN(n2281) );
  NOR2_X1 U1980 ( .A1(n974), .A2(n2258), .ZN(n1857) );
  OAI22_X1 U1981 ( .A1(n878), .A2(n2275), .B1(n334), .B2(n2256), .ZN(n1856) );
  OAI22_X1 U1982 ( .A1(n78), .A2(n2251), .B1(n526), .B2(n2253), .ZN(n1855) );
  OAI22_X1 U1983 ( .A1(n686), .A2(n2262), .B1(n782), .B2(n2279), .ZN(n1854) );
  NOR4_X1 U1984 ( .A1(n1857), .A2(n1856), .A3(n1855), .A4(n1854), .ZN(n1873)
         );
  OAI22_X1 U1985 ( .A1(n622), .A2(n1678), .B1(n110), .B2(n2274), .ZN(n1861) );
  OAI22_X1 U1986 ( .A1(n462), .A2(n2268), .B1(n942), .B2(n2277), .ZN(n1860) );
  OAI22_X1 U1987 ( .A1(n750), .A2(n2276), .B1(n846), .B2(n2261), .ZN(n1859) );
  OAI22_X1 U1988 ( .A1(n366), .A2(n2260), .B1(n558), .B2(n2265), .ZN(n1858) );
  NOR4_X1 U1989 ( .A1(n1861), .A2(n1860), .A3(n1859), .A4(n1858), .ZN(n1872)
         );
  OAI22_X1 U1990 ( .A1(n14), .A2(n2264), .B1(n718), .B2(n2269), .ZN(n1865) );
  OAI22_X1 U1991 ( .A1(n910), .A2(n2272), .B1(n398), .B2(n2270), .ZN(n1864) );
  OAI22_X1 U1992 ( .A1(n654), .A2(n2278), .B1(n814), .B2(n2273), .ZN(n1863) );
  OAI22_X1 U1993 ( .A1(n206), .A2(n2266), .B1(n302), .B2(n2280), .ZN(n1862) );
  NOR4_X1 U1994 ( .A1(n1865), .A2(n1864), .A3(n1863), .A4(n1862), .ZN(n1871)
         );
  OAI22_X1 U1995 ( .A1(n494), .A2(n2259), .B1(n46), .B2(n2255), .ZN(n1869) );
  OAI22_X1 U1996 ( .A1(n590), .A2(n2250), .B1(n270), .B2(n2252), .ZN(n1868) );
  OAI22_X1 U1997 ( .A1(n430), .A2(n2267), .B1(n142), .B2(n2254), .ZN(n1867) );
  OAI22_X1 U1998 ( .A1(n238), .A2(n2263), .B1(n174), .B2(n2257), .ZN(n1866) );
  NOR4_X1 U1999 ( .A1(n1869), .A2(n1868), .A3(n1867), .A4(n1866), .ZN(n1870)
         );
  NAND4_X1 U2000 ( .A1(n1873), .A2(n1872), .A3(n1871), .A4(n1870), .ZN(n1874)
         );
  AOI22_X1 U2001 ( .A1(n1680), .A2(n1874), .B1(n1679), .B2(lo_out[13]), .ZN(
        n1875) );
  OAI21_X1 U2002 ( .B1(n2283), .B2(n1632), .A(n1875), .ZN(rp1[13]) );
  NOR2_X1 U2003 ( .A1(n367), .A2(n2260), .ZN(n1879) );
  OAI22_X1 U2004 ( .A1(n143), .A2(n2254), .B1(n911), .B2(n2272), .ZN(n1878) );
  OAI22_X1 U2005 ( .A1(n591), .A2(n2250), .B1(n815), .B2(n2273), .ZN(n1877) );
  OAI22_X1 U2006 ( .A1(n527), .A2(n2253), .B1(n47), .B2(n2255), .ZN(n1876) );
  NOR4_X1 U2007 ( .A1(n1879), .A2(n1878), .A3(n1877), .A4(n1876), .ZN(n1895)
         );
  OAI22_X1 U2008 ( .A1(n943), .A2(n2277), .B1(n335), .B2(n2256), .ZN(n1883) );
  OAI22_X1 U2009 ( .A1(n687), .A2(n2262), .B1(n655), .B2(n2278), .ZN(n1882) );
  OAI22_X1 U2010 ( .A1(n879), .A2(n2275), .B1(n271), .B2(n2252), .ZN(n1881) );
  OAI22_X1 U2011 ( .A1(n783), .A2(n2279), .B1(n559), .B2(n2265), .ZN(n1880) );
  NOR4_X1 U2012 ( .A1(n1883), .A2(n1882), .A3(n1881), .A4(n1880), .ZN(n1894)
         );
  OAI22_X1 U2013 ( .A1(n175), .A2(n2257), .B1(n15), .B2(n2264), .ZN(n1887) );
  OAI22_X1 U2014 ( .A1(n303), .A2(n2280), .B1(n719), .B2(n2269), .ZN(n1886) );
  OAI22_X1 U2015 ( .A1(n79), .A2(n2251), .B1(n847), .B2(n2261), .ZN(n1885) );
  OAI22_X1 U2016 ( .A1(n399), .A2(n2270), .B1(n431), .B2(n2267), .ZN(n1884) );
  NOR4_X1 U2017 ( .A1(n1887), .A2(n1886), .A3(n1885), .A4(n1884), .ZN(n1893)
         );
  OAI22_X1 U2018 ( .A1(n751), .A2(n2276), .B1(n623), .B2(n2271), .ZN(n1891) );
  OAI22_X1 U2019 ( .A1(n111), .A2(n2274), .B1(n495), .B2(n2259), .ZN(n1890) );
  OAI22_X1 U2020 ( .A1(n207), .A2(n2266), .B1(n975), .B2(n2258), .ZN(n1889) );
  OAI22_X1 U2021 ( .A1(n239), .A2(n2263), .B1(n463), .B2(n2268), .ZN(n1888) );
  NOR4_X1 U2022 ( .A1(n1891), .A2(n1890), .A3(n1889), .A4(n1888), .ZN(n1892)
         );
  NAND4_X1 U2023 ( .A1(n1895), .A2(n1894), .A3(n1893), .A4(n1892), .ZN(n1896)
         );
  AOI22_X1 U2024 ( .A1(n1680), .A2(n1896), .B1(n1679), .B2(lo_out[14]), .ZN(
        n1897) );
  OAI21_X1 U2025 ( .B1(n2283), .B2(n1633), .A(n1897), .ZN(rp1[14]) );
  NOR2_X1 U2026 ( .A1(n496), .A2(n2259), .ZN(n1901) );
  OAI22_X1 U2027 ( .A1(n656), .A2(n2278), .B1(n176), .B2(n2257), .ZN(n1900) );
  OAI22_X1 U2028 ( .A1(n592), .A2(n2250), .B1(n688), .B2(n2262), .ZN(n1899) );
  OAI22_X1 U2029 ( .A1(n336), .A2(n2256), .B1(n848), .B2(n2261), .ZN(n1898) );
  NOR4_X1 U2030 ( .A1(n1901), .A2(n1900), .A3(n1899), .A4(n1898), .ZN(n1917)
         );
  OAI22_X1 U2031 ( .A1(n272), .A2(n2252), .B1(n816), .B2(n2273), .ZN(n1905) );
  OAI22_X1 U2032 ( .A1(n752), .A2(n2276), .B1(n624), .B2(n2271), .ZN(n1904) );
  OAI22_X1 U2033 ( .A1(n16), .A2(n2264), .B1(n304), .B2(n2280), .ZN(n1903) );
  OAI22_X1 U2034 ( .A1(n464), .A2(n2268), .B1(n144), .B2(n2254), .ZN(n1902) );
  NOR4_X1 U2035 ( .A1(n1905), .A2(n1904), .A3(n1903), .A4(n1902), .ZN(n1916)
         );
  OAI22_X1 U2036 ( .A1(n912), .A2(n2272), .B1(n112), .B2(n2274), .ZN(n1909) );
  OAI22_X1 U2037 ( .A1(n400), .A2(n2270), .B1(n80), .B2(n2251), .ZN(n1908) );
  OAI22_X1 U2038 ( .A1(n528), .A2(n2253), .B1(n240), .B2(n2263), .ZN(n1907) );
  OAI22_X1 U2039 ( .A1(n208), .A2(n2266), .B1(n944), .B2(n2277), .ZN(n1906) );
  NOR4_X1 U2040 ( .A1(n1909), .A2(n1908), .A3(n1907), .A4(n1906), .ZN(n1915)
         );
  OAI22_X1 U2041 ( .A1(n784), .A2(n2279), .B1(n880), .B2(n2275), .ZN(n1913) );
  OAI22_X1 U2042 ( .A1(n560), .A2(n2265), .B1(n432), .B2(n2267), .ZN(n1912) );
  OAI22_X1 U2043 ( .A1(n976), .A2(n2258), .B1(n48), .B2(n2255), .ZN(n1911) );
  OAI22_X1 U2044 ( .A1(n720), .A2(n2269), .B1(n368), .B2(n2260), .ZN(n1910) );
  NOR4_X1 U2045 ( .A1(n1913), .A2(n1912), .A3(n1911), .A4(n1910), .ZN(n1914)
         );
  NAND4_X1 U2046 ( .A1(n1917), .A2(n1916), .A3(n1915), .A4(n1914), .ZN(n1918)
         );
  AOI22_X1 U2047 ( .A1(n2282), .A2(n1918), .B1(n1679), .B2(lo_out[15]), .ZN(
        n1919) );
  OAI21_X1 U2048 ( .B1(n2283), .B2(n1634), .A(n1919), .ZN(rp1[15]) );
  NOR2_X1 U2049 ( .A1(n593), .A2(n2250), .ZN(n1923) );
  OAI22_X1 U2050 ( .A1(n49), .A2(n2255), .B1(n913), .B2(n2272), .ZN(n1922) );
  OAI22_X1 U2051 ( .A1(n241), .A2(n2263), .B1(n689), .B2(n2262), .ZN(n1921) );
  OAI22_X1 U2052 ( .A1(n497), .A2(n2259), .B1(n273), .B2(n2252), .ZN(n1920) );
  NOR4_X1 U2053 ( .A1(n1923), .A2(n1922), .A3(n1921), .A4(n1920), .ZN(n1939)
         );
  OAI22_X1 U2054 ( .A1(n817), .A2(n2273), .B1(n401), .B2(n2270), .ZN(n1927) );
  OAI22_X1 U2055 ( .A1(n465), .A2(n2268), .B1(n305), .B2(n2280), .ZN(n1926) );
  OAI22_X1 U2056 ( .A1(n145), .A2(n2254), .B1(n113), .B2(n2274), .ZN(n1925) );
  OAI22_X1 U2057 ( .A1(n369), .A2(n2260), .B1(n177), .B2(n2257), .ZN(n1924) );
  NOR4_X1 U2058 ( .A1(n1927), .A2(n1926), .A3(n1925), .A4(n1924), .ZN(n1938)
         );
  OAI22_X1 U2059 ( .A1(n945), .A2(n2277), .B1(n529), .B2(n2253), .ZN(n1931) );
  OAI22_X1 U2060 ( .A1(n17), .A2(n2264), .B1(n625), .B2(n2271), .ZN(n1930) );
  OAI22_X1 U2061 ( .A1(n753), .A2(n2276), .B1(n849), .B2(n2261), .ZN(n1929) );
  OAI22_X1 U2062 ( .A1(n881), .A2(n2275), .B1(n337), .B2(n2256), .ZN(n1928) );
  NOR4_X1 U2063 ( .A1(n1931), .A2(n1930), .A3(n1929), .A4(n1928), .ZN(n1937)
         );
  OAI22_X1 U2064 ( .A1(n785), .A2(n2279), .B1(n209), .B2(n2266), .ZN(n1935) );
  OAI22_X1 U2065 ( .A1(n721), .A2(n2269), .B1(n657), .B2(n2278), .ZN(n1934) );
  OAI22_X1 U2066 ( .A1(n561), .A2(n2265), .B1(n977), .B2(n2258), .ZN(n1933) );
  OAI22_X1 U2067 ( .A1(n433), .A2(n2267), .B1(n81), .B2(n2251), .ZN(n1932) );
  NOR4_X1 U2068 ( .A1(n1935), .A2(n1934), .A3(n1933), .A4(n1932), .ZN(n1936)
         );
  NAND4_X1 U2069 ( .A1(n1939), .A2(n1938), .A3(n1937), .A4(n1936), .ZN(n1940)
         );
  AOI22_X1 U2070 ( .A1(n2282), .A2(n1940), .B1(n2281), .B2(lo_out[16]), .ZN(
        n1941) );
  OAI21_X1 U2071 ( .B1(n2283), .B2(n1635), .A(n1941), .ZN(rp1[16]) );
  NOR2_X1 U2072 ( .A1(n178), .A2(n2257), .ZN(n1945) );
  OAI22_X1 U2073 ( .A1(n306), .A2(n2280), .B1(n18), .B2(n2264), .ZN(n1944) );
  OAI22_X1 U2074 ( .A1(n242), .A2(n2263), .B1(n466), .B2(n2268), .ZN(n1943) );
  OAI22_X1 U2075 ( .A1(n434), .A2(n2267), .B1(n946), .B2(n2277), .ZN(n1942) );
  NOR4_X1 U2076 ( .A1(n1945), .A2(n1944), .A3(n1943), .A4(n1942), .ZN(n1961)
         );
  OAI22_X1 U2077 ( .A1(n786), .A2(n2279), .B1(n498), .B2(n2259), .ZN(n1949) );
  OAI22_X1 U2078 ( .A1(n530), .A2(n2253), .B1(n370), .B2(n2260), .ZN(n1948) );
  OAI22_X1 U2079 ( .A1(n338), .A2(n2256), .B1(n562), .B2(n2265), .ZN(n1947) );
  OAI22_X1 U2080 ( .A1(n50), .A2(n2255), .B1(n658), .B2(n2278), .ZN(n1946) );
  NOR4_X1 U2081 ( .A1(n1949), .A2(n1948), .A3(n1947), .A4(n1946), .ZN(n1960)
         );
  OAI22_X1 U2082 ( .A1(n722), .A2(n2269), .B1(n882), .B2(n2275), .ZN(n1953) );
  OAI22_X1 U2083 ( .A1(n850), .A2(n2261), .B1(n626), .B2(n2271), .ZN(n1952) );
  OAI22_X1 U2084 ( .A1(n402), .A2(n2270), .B1(n594), .B2(n2250), .ZN(n1951) );
  OAI22_X1 U2085 ( .A1(n274), .A2(n2252), .B1(n114), .B2(n2274), .ZN(n1950) );
  NOR4_X1 U2086 ( .A1(n1953), .A2(n1952), .A3(n1951), .A4(n1950), .ZN(n1959)
         );
  OAI22_X1 U2087 ( .A1(n82), .A2(n2251), .B1(n818), .B2(n2273), .ZN(n1957) );
  OAI22_X1 U2088 ( .A1(n914), .A2(n2272), .B1(n690), .B2(n2262), .ZN(n1956) );
  OAI22_X1 U2089 ( .A1(n978), .A2(n2258), .B1(n210), .B2(n2266), .ZN(n1955) );
  OAI22_X1 U2090 ( .A1(n754), .A2(n2276), .B1(n146), .B2(n2254), .ZN(n1954) );
  NOR4_X1 U2091 ( .A1(n1957), .A2(n1956), .A3(n1955), .A4(n1954), .ZN(n1958)
         );
  NAND4_X1 U2092 ( .A1(n1961), .A2(n1960), .A3(n1959), .A4(n1958), .ZN(n1962)
         );
  AOI22_X1 U2093 ( .A1(n2282), .A2(n1962), .B1(n1679), .B2(lo_out[17]), .ZN(
        n1963) );
  OAI21_X1 U2094 ( .B1(n2283), .B2(n1650), .A(n1963), .ZN(rp1[17]) );
  NOR2_X1 U2095 ( .A1(n947), .A2(n2277), .ZN(n1967) );
  OAI22_X1 U2096 ( .A1(n211), .A2(n2266), .B1(n307), .B2(n2280), .ZN(n1966) );
  OAI22_X1 U2097 ( .A1(n627), .A2(n2271), .B1(n755), .B2(n2276), .ZN(n1965) );
  OAI22_X1 U2098 ( .A1(n819), .A2(n2273), .B1(n787), .B2(n2279), .ZN(n1964) );
  NOR4_X1 U2099 ( .A1(n1967), .A2(n1966), .A3(n1965), .A4(n1964), .ZN(n1983)
         );
  OAI22_X1 U2100 ( .A1(n19), .A2(n2264), .B1(n371), .B2(n2260), .ZN(n1971) );
  OAI22_X1 U2101 ( .A1(n435), .A2(n2267), .B1(n915), .B2(n2272), .ZN(n1970) );
  OAI22_X1 U2102 ( .A1(n659), .A2(n2278), .B1(n499), .B2(n2259), .ZN(n1969) );
  OAI22_X1 U2103 ( .A1(n531), .A2(n2253), .B1(n563), .B2(n2265), .ZN(n1968) );
  NOR4_X1 U2104 ( .A1(n1971), .A2(n1970), .A3(n1969), .A4(n1968), .ZN(n1982)
         );
  OAI22_X1 U2105 ( .A1(n83), .A2(n2251), .B1(n243), .B2(n2263), .ZN(n1975) );
  OAI22_X1 U2106 ( .A1(n403), .A2(n2270), .B1(n147), .B2(n2254), .ZN(n1974) );
  OAI22_X1 U2107 ( .A1(n723), .A2(n2269), .B1(n979), .B2(n2258), .ZN(n1973) );
  OAI22_X1 U2108 ( .A1(n51), .A2(n2255), .B1(n691), .B2(n2262), .ZN(n1972) );
  NOR4_X1 U2109 ( .A1(n1975), .A2(n1974), .A3(n1973), .A4(n1972), .ZN(n1981)
         );
  OAI22_X1 U2110 ( .A1(n275), .A2(n2252), .B1(n467), .B2(n2268), .ZN(n1979) );
  OAI22_X1 U2111 ( .A1(n339), .A2(n2256), .B1(n179), .B2(n2257), .ZN(n1978) );
  OAI22_X1 U2112 ( .A1(n595), .A2(n2250), .B1(n115), .B2(n2274), .ZN(n1977) );
  OAI22_X1 U2113 ( .A1(n851), .A2(n2261), .B1(n883), .B2(n2275), .ZN(n1976) );
  NOR4_X1 U2114 ( .A1(n1979), .A2(n1978), .A3(n1977), .A4(n1976), .ZN(n1980)
         );
  NAND4_X1 U2115 ( .A1(n1983), .A2(n1982), .A3(n1981), .A4(n1980), .ZN(n1984)
         );
  AOI22_X1 U2116 ( .A1(n2282), .A2(n1984), .B1(n2281), .B2(lo_out[18]), .ZN(
        n1985) );
  OAI21_X1 U2117 ( .B1(n2283), .B2(n1636), .A(n1985), .ZN(rp1[18]) );
  NOR2_X1 U2118 ( .A1(n696), .A2(n2262), .ZN(n1989) );
  OAI22_X1 U2119 ( .A1(n536), .A2(n2253), .B1(n88), .B2(n2251), .ZN(n1988) );
  OAI22_X1 U2120 ( .A1(n664), .A2(n2278), .B1(n504), .B2(n2259), .ZN(n1987) );
  OAI22_X1 U2121 ( .A1(n568), .A2(n2265), .B1(n472), .B2(n2268), .ZN(n1986) );
  NOR4_X1 U2122 ( .A1(n1989), .A2(n1988), .A3(n1987), .A4(n1986), .ZN(n2005)
         );
  OAI22_X1 U2123 ( .A1(n760), .A2(n2276), .B1(n984), .B2(n2258), .ZN(n1993) );
  OAI22_X1 U2124 ( .A1(n248), .A2(n2263), .B1(n728), .B2(n2269), .ZN(n1992) );
  OAI22_X1 U2125 ( .A1(n888), .A2(n2275), .B1(n312), .B2(n2280), .ZN(n1991) );
  OAI22_X1 U2126 ( .A1(n152), .A2(n1677), .B1(n24), .B2(n2264), .ZN(n1990) );
  NOR4_X1 U2127 ( .A1(n1993), .A2(n1992), .A3(n1991), .A4(n1990), .ZN(n2004)
         );
  OAI22_X1 U2128 ( .A1(n600), .A2(n2250), .B1(n408), .B2(n2270), .ZN(n1997) );
  OAI22_X1 U2129 ( .A1(n280), .A2(n2252), .B1(n376), .B2(n2260), .ZN(n1996) );
  OAI22_X1 U2130 ( .A1(n184), .A2(n2257), .B1(n952), .B2(n2277), .ZN(n1995) );
  OAI22_X1 U2131 ( .A1(n792), .A2(n2279), .B1(n344), .B2(n2256), .ZN(n1994) );
  NOR4_X1 U2132 ( .A1(n1997), .A2(n1996), .A3(n1995), .A4(n1994), .ZN(n2003)
         );
  OAI22_X1 U2133 ( .A1(n856), .A2(n2261), .B1(n216), .B2(n2266), .ZN(n2001) );
  OAI22_X1 U2134 ( .A1(n56), .A2(n2255), .B1(n632), .B2(n2271), .ZN(n2000) );
  OAI22_X1 U2135 ( .A1(n440), .A2(n2267), .B1(n120), .B2(n2274), .ZN(n1999) );
  OAI22_X1 U2136 ( .A1(n920), .A2(n2272), .B1(n824), .B2(n2273), .ZN(n1998) );
  NOR4_X1 U2137 ( .A1(n2001), .A2(n2000), .A3(n1999), .A4(n1998), .ZN(n2002)
         );
  NAND4_X1 U2138 ( .A1(n2005), .A2(n2004), .A3(n2003), .A4(n2002), .ZN(n2006)
         );
  AOI22_X1 U2139 ( .A1(n1680), .A2(n2006), .B1(n2281), .B2(lo_out[23]), .ZN(
        n2007) );
  OAI21_X1 U2140 ( .B1(n2283), .B2(n1641), .A(n2007), .ZN(rp1[23]) );
  NOR2_X1 U2141 ( .A1(n633), .A2(n2271), .ZN(n2011) );
  OAI22_X1 U2142 ( .A1(n921), .A2(n2272), .B1(n153), .B2(n2254), .ZN(n2010) );
  OAI22_X1 U2143 ( .A1(n537), .A2(n2253), .B1(n665), .B2(n2278), .ZN(n2009) );
  OAI22_X1 U2144 ( .A1(n313), .A2(n2280), .B1(n121), .B2(n2274), .ZN(n2008) );
  NOR4_X1 U2145 ( .A1(n2011), .A2(n2010), .A3(n2009), .A4(n2008), .ZN(n2027)
         );
  OAI22_X1 U2146 ( .A1(n345), .A2(n2256), .B1(n409), .B2(n2270), .ZN(n2015) );
  OAI22_X1 U2147 ( .A1(n441), .A2(n2267), .B1(n889), .B2(n2275), .ZN(n2014) );
  OAI22_X1 U2148 ( .A1(n473), .A2(n2268), .B1(n25), .B2(n2264), .ZN(n2013) );
  OAI22_X1 U2149 ( .A1(n569), .A2(n2265), .B1(n793), .B2(n2279), .ZN(n2012) );
  NOR4_X1 U2150 ( .A1(n2015), .A2(n2014), .A3(n2013), .A4(n2012), .ZN(n2026)
         );
  OAI22_X1 U2151 ( .A1(n825), .A2(n2273), .B1(n505), .B2(n2259), .ZN(n2019) );
  OAI22_X1 U2152 ( .A1(n601), .A2(n2250), .B1(n249), .B2(n2263), .ZN(n2018) );
  OAI22_X1 U2153 ( .A1(n985), .A2(n2258), .B1(n697), .B2(n2262), .ZN(n2017) );
  OAI22_X1 U2154 ( .A1(n281), .A2(n2252), .B1(n729), .B2(n2269), .ZN(n2016) );
  NOR4_X1 U2155 ( .A1(n2019), .A2(n2018), .A3(n2017), .A4(n2016), .ZN(n2025)
         );
  OAI22_X1 U2156 ( .A1(n185), .A2(n2257), .B1(n57), .B2(n2255), .ZN(n2023) );
  OAI22_X1 U2157 ( .A1(n953), .A2(n2277), .B1(n857), .B2(n2261), .ZN(n2022) );
  OAI22_X1 U2158 ( .A1(n217), .A2(n2266), .B1(n89), .B2(n2251), .ZN(n2021) );
  OAI22_X1 U2159 ( .A1(n761), .A2(n2276), .B1(n377), .B2(n2260), .ZN(n2020) );
  NOR4_X1 U2160 ( .A1(n2023), .A2(n2022), .A3(n2021), .A4(n2020), .ZN(n2024)
         );
  NAND4_X1 U2161 ( .A1(n2027), .A2(n2026), .A3(n2025), .A4(n2024), .ZN(n2028)
         );
  AOI22_X1 U2162 ( .A1(n1680), .A2(n2028), .B1(n2281), .B2(lo_out[24]), .ZN(
        n2029) );
  OAI21_X1 U2163 ( .B1(n2283), .B2(n1642), .A(n2029), .ZN(rp1[24]) );
  NOR2_X1 U2164 ( .A1(n186), .A2(n2257), .ZN(n2033) );
  OAI22_X1 U2165 ( .A1(n890), .A2(n2275), .B1(n378), .B2(n2260), .ZN(n2032) );
  OAI22_X1 U2166 ( .A1(n762), .A2(n2276), .B1(n826), .B2(n2273), .ZN(n2031) );
  OAI22_X1 U2167 ( .A1(n538), .A2(n2253), .B1(n58), .B2(n2255), .ZN(n2030) );
  NOR4_X1 U2168 ( .A1(n2033), .A2(n2032), .A3(n2031), .A4(n2030), .ZN(n2049)
         );
  OAI22_X1 U2169 ( .A1(n442), .A2(n2267), .B1(n410), .B2(n2270), .ZN(n2037) );
  OAI22_X1 U2170 ( .A1(n282), .A2(n2252), .B1(n26), .B2(n2264), .ZN(n2036) );
  OAI22_X1 U2171 ( .A1(n122), .A2(n2274), .B1(n730), .B2(n2269), .ZN(n2035) );
  OAI22_X1 U2172 ( .A1(n90), .A2(n2251), .B1(n154), .B2(n1677), .ZN(n2034) );
  NOR4_X1 U2173 ( .A1(n2037), .A2(n2036), .A3(n2035), .A4(n2034), .ZN(n2048)
         );
  OAI22_X1 U2174 ( .A1(n250), .A2(n2263), .B1(n474), .B2(n2268), .ZN(n2041) );
  OAI22_X1 U2175 ( .A1(n922), .A2(n2272), .B1(n570), .B2(n2265), .ZN(n2040) );
  OAI22_X1 U2176 ( .A1(n858), .A2(n2261), .B1(n666), .B2(n2278), .ZN(n2039) );
  OAI22_X1 U2177 ( .A1(n602), .A2(n2250), .B1(n986), .B2(n2258), .ZN(n2038) );
  NOR4_X1 U2178 ( .A1(n2041), .A2(n2040), .A3(n2039), .A4(n2038), .ZN(n2047)
         );
  OAI22_X1 U2179 ( .A1(n954), .A2(n2277), .B1(n698), .B2(n2262), .ZN(n2045) );
  OAI22_X1 U2180 ( .A1(n346), .A2(n2256), .B1(n218), .B2(n2266), .ZN(n2044) );
  OAI22_X1 U2181 ( .A1(n634), .A2(n2271), .B1(n506), .B2(n2259), .ZN(n2043) );
  OAI22_X1 U2182 ( .A1(n794), .A2(n2279), .B1(n314), .B2(n2280), .ZN(n2042) );
  NOR4_X1 U2183 ( .A1(n2045), .A2(n2044), .A3(n2043), .A4(n2042), .ZN(n2046)
         );
  NAND4_X1 U2184 ( .A1(n2049), .A2(n2048), .A3(n2047), .A4(n2046), .ZN(n2050)
         );
  AOI22_X1 U2185 ( .A1(n2282), .A2(n2050), .B1(n1679), .B2(lo_out[25]), .ZN(
        n2051) );
  OAI21_X1 U2186 ( .B1(n2283), .B2(n1652), .A(n2051), .ZN(rp1[25]) );
  NOR2_X1 U2187 ( .A1(n955), .A2(n2277), .ZN(n2055) );
  OAI22_X1 U2188 ( .A1(n763), .A2(n2276), .B1(n923), .B2(n2272), .ZN(n2054) );
  OAI22_X1 U2189 ( .A1(n635), .A2(n2271), .B1(n379), .B2(n2260), .ZN(n2053) );
  OAI22_X1 U2190 ( .A1(n315), .A2(n2280), .B1(n251), .B2(n2263), .ZN(n2052) );
  NOR4_X1 U2191 ( .A1(n2055), .A2(n2054), .A3(n2053), .A4(n2052), .ZN(n2071)
         );
  OAI22_X1 U2192 ( .A1(n731), .A2(n2269), .B1(n539), .B2(n2253), .ZN(n2059) );
  OAI22_X1 U2193 ( .A1(n827), .A2(n2273), .B1(n347), .B2(n2256), .ZN(n2058) );
  OAI22_X1 U2194 ( .A1(n475), .A2(n2268), .B1(n59), .B2(n2255), .ZN(n2057) );
  OAI22_X1 U2195 ( .A1(n443), .A2(n2267), .B1(n91), .B2(n2251), .ZN(n2056) );
  NOR4_X1 U2196 ( .A1(n2059), .A2(n2058), .A3(n2057), .A4(n2056), .ZN(n2070)
         );
  OAI22_X1 U2197 ( .A1(n891), .A2(n2275), .B1(n987), .B2(n2258), .ZN(n2063) );
  OAI22_X1 U2198 ( .A1(n123), .A2(n2274), .B1(n187), .B2(n2257), .ZN(n2062) );
  OAI22_X1 U2199 ( .A1(n859), .A2(n2261), .B1(n795), .B2(n2279), .ZN(n2061) );
  OAI22_X1 U2200 ( .A1(n411), .A2(n2270), .B1(n699), .B2(n2262), .ZN(n2060) );
  NOR4_X1 U2201 ( .A1(n2063), .A2(n2062), .A3(n2061), .A4(n2060), .ZN(n2069)
         );
  OAI22_X1 U2202 ( .A1(n283), .A2(n2252), .B1(n603), .B2(n2250), .ZN(n2067) );
  OAI22_X1 U2203 ( .A1(n507), .A2(n2259), .B1(n571), .B2(n2265), .ZN(n2066) );
  OAI22_X1 U2204 ( .A1(n27), .A2(n2264), .B1(n155), .B2(n1677), .ZN(n2065) );
  OAI22_X1 U2205 ( .A1(n219), .A2(n2266), .B1(n667), .B2(n2278), .ZN(n2064) );
  NOR4_X1 U2206 ( .A1(n2067), .A2(n2066), .A3(n2065), .A4(n2064), .ZN(n2068)
         );
  NAND4_X1 U2207 ( .A1(n2071), .A2(n2070), .A3(n2069), .A4(n2068), .ZN(n2072)
         );
  AOI22_X1 U2208 ( .A1(n1680), .A2(n2072), .B1(n1679), .B2(lo_out[26]), .ZN(
        n2073) );
  OAI21_X1 U2209 ( .B1(n2283), .B2(n1643), .A(n2073), .ZN(rp1[26]) );
  NOR2_X1 U2210 ( .A1(n156), .A2(n2254), .ZN(n2077) );
  OAI22_X1 U2211 ( .A1(n860), .A2(n2261), .B1(n252), .B2(n2263), .ZN(n2076) );
  OAI22_X1 U2212 ( .A1(n732), .A2(n2269), .B1(n924), .B2(n2272), .ZN(n2075) );
  OAI22_X1 U2213 ( .A1(n220), .A2(n2266), .B1(n124), .B2(n2274), .ZN(n2074) );
  NOR4_X1 U2214 ( .A1(n2077), .A2(n2076), .A3(n2075), .A4(n2074), .ZN(n2093)
         );
  OAI22_X1 U2215 ( .A1(n348), .A2(n2256), .B1(n284), .B2(n2252), .ZN(n2081) );
  OAI22_X1 U2216 ( .A1(n60), .A2(n2255), .B1(n444), .B2(n2267), .ZN(n2080) );
  OAI22_X1 U2217 ( .A1(n188), .A2(n2257), .B1(n796), .B2(n2279), .ZN(n2079) );
  OAI22_X1 U2218 ( .A1(n508), .A2(n2259), .B1(n604), .B2(n2250), .ZN(n2078) );
  NOR4_X1 U2219 ( .A1(n2081), .A2(n2080), .A3(n2079), .A4(n2078), .ZN(n2092)
         );
  OAI22_X1 U2220 ( .A1(n28), .A2(n2264), .B1(n476), .B2(n2268), .ZN(n2085) );
  OAI22_X1 U2221 ( .A1(n540), .A2(n2253), .B1(n412), .B2(n2270), .ZN(n2084) );
  OAI22_X1 U2222 ( .A1(n828), .A2(n2273), .B1(n92), .B2(n2251), .ZN(n2083) );
  OAI22_X1 U2223 ( .A1(n892), .A2(n2275), .B1(n764), .B2(n2276), .ZN(n2082) );
  NOR4_X1 U2224 ( .A1(n2085), .A2(n2084), .A3(n2083), .A4(n2082), .ZN(n2091)
         );
  OAI22_X1 U2225 ( .A1(n380), .A2(n2260), .B1(n572), .B2(n2265), .ZN(n2089) );
  OAI22_X1 U2226 ( .A1(n668), .A2(n2278), .B1(n988), .B2(n2258), .ZN(n2088) );
  OAI22_X1 U2227 ( .A1(n956), .A2(n2277), .B1(n636), .B2(n1678), .ZN(n2087) );
  OAI22_X1 U2228 ( .A1(n316), .A2(n2280), .B1(n700), .B2(n2262), .ZN(n2086) );
  NOR4_X1 U2229 ( .A1(n2089), .A2(n2088), .A3(n2087), .A4(n2086), .ZN(n2090)
         );
  NAND4_X1 U2230 ( .A1(n2093), .A2(n2092), .A3(n2091), .A4(n2090), .ZN(n2094)
         );
  AOI22_X1 U2231 ( .A1(n1680), .A2(n2094), .B1(n2281), .B2(lo_out[27]), .ZN(
        n2095) );
  OAI21_X1 U2232 ( .B1(n2283), .B2(n1644), .A(n2095), .ZN(rp1[27]) );
  NOR2_X1 U2233 ( .A1(n573), .A2(n2265), .ZN(n2099) );
  OAI22_X1 U2234 ( .A1(n317), .A2(n2280), .B1(n285), .B2(n2252), .ZN(n2098) );
  OAI22_X1 U2235 ( .A1(n701), .A2(n2262), .B1(n669), .B2(n2278), .ZN(n2097) );
  OAI22_X1 U2236 ( .A1(n509), .A2(n2259), .B1(n765), .B2(n2276), .ZN(n2096) );
  NOR4_X1 U2237 ( .A1(n2099), .A2(n2098), .A3(n2097), .A4(n2096), .ZN(n2115)
         );
  OAI22_X1 U2238 ( .A1(n93), .A2(n2251), .B1(n893), .B2(n2275), .ZN(n2103) );
  OAI22_X1 U2239 ( .A1(n477), .A2(n2268), .B1(n541), .B2(n2253), .ZN(n2102) );
  OAI22_X1 U2240 ( .A1(n221), .A2(n2266), .B1(n829), .B2(n2273), .ZN(n2101) );
  OAI22_X1 U2241 ( .A1(n797), .A2(n2279), .B1(n349), .B2(n2256), .ZN(n2100) );
  NOR4_X1 U2242 ( .A1(n2103), .A2(n2102), .A3(n2101), .A4(n2100), .ZN(n2114)
         );
  OAI22_X1 U2243 ( .A1(n157), .A2(n1677), .B1(n733), .B2(n2269), .ZN(n2107) );
  OAI22_X1 U2244 ( .A1(n605), .A2(n2250), .B1(n925), .B2(n2272), .ZN(n2106) );
  OAI22_X1 U2245 ( .A1(n637), .A2(n2271), .B1(n989), .B2(n2258), .ZN(n2105) );
  OAI22_X1 U2246 ( .A1(n957), .A2(n2277), .B1(n413), .B2(n2270), .ZN(n2104) );
  NOR4_X1 U2247 ( .A1(n2107), .A2(n2106), .A3(n2105), .A4(n2104), .ZN(n2113)
         );
  OAI22_X1 U2248 ( .A1(n253), .A2(n2263), .B1(n29), .B2(n2264), .ZN(n2111) );
  OAI22_X1 U2249 ( .A1(n189), .A2(n2257), .B1(n861), .B2(n2261), .ZN(n2110) );
  OAI22_X1 U2250 ( .A1(n125), .A2(n2274), .B1(n61), .B2(n2255), .ZN(n2109) );
  OAI22_X1 U2251 ( .A1(n445), .A2(n2267), .B1(n381), .B2(n2260), .ZN(n2108) );
  NOR4_X1 U2252 ( .A1(n2111), .A2(n2110), .A3(n2109), .A4(n2108), .ZN(n2112)
         );
  NAND4_X1 U2253 ( .A1(n2115), .A2(n2114), .A3(n2113), .A4(n2112), .ZN(n2116)
         );
  AOI22_X1 U2254 ( .A1(n1680), .A2(n2116), .B1(n2281), .B2(lo_out[28]), .ZN(
        n2117) );
  OAI21_X1 U2255 ( .B1(n2283), .B2(n1645), .A(n2117), .ZN(rp1[28]) );
  NOR2_X1 U2256 ( .A1(n94), .A2(n2251), .ZN(n2121) );
  OAI22_X1 U2257 ( .A1(n830), .A2(n2273), .B1(n734), .B2(n2269), .ZN(n2120) );
  OAI22_X1 U2258 ( .A1(n478), .A2(n2268), .B1(n350), .B2(n2256), .ZN(n2119) );
  OAI22_X1 U2259 ( .A1(n318), .A2(n2280), .B1(n222), .B2(n2266), .ZN(n2118) );
  NOR4_X1 U2260 ( .A1(n2121), .A2(n2120), .A3(n2119), .A4(n2118), .ZN(n2137)
         );
  OAI22_X1 U2261 ( .A1(n958), .A2(n2277), .B1(n638), .B2(n2271), .ZN(n2125) );
  OAI22_X1 U2262 ( .A1(n126), .A2(n2274), .B1(n542), .B2(n2253), .ZN(n2124) );
  OAI22_X1 U2263 ( .A1(n446), .A2(n2267), .B1(n30), .B2(n2264), .ZN(n2123) );
  OAI22_X1 U2264 ( .A1(n894), .A2(n2275), .B1(n510), .B2(n2259), .ZN(n2122) );
  NOR4_X1 U2265 ( .A1(n2125), .A2(n2124), .A3(n2123), .A4(n2122), .ZN(n2136)
         );
  OAI22_X1 U2266 ( .A1(n62), .A2(n2255), .B1(n798), .B2(n2279), .ZN(n2129) );
  OAI22_X1 U2267 ( .A1(n670), .A2(n2278), .B1(n382), .B2(n2260), .ZN(n2128) );
  OAI22_X1 U2268 ( .A1(n926), .A2(n2272), .B1(n862), .B2(n2261), .ZN(n2127) );
  OAI22_X1 U2269 ( .A1(n190), .A2(n2257), .B1(n158), .B2(n1677), .ZN(n2126) );
  NOR4_X1 U2270 ( .A1(n2129), .A2(n2128), .A3(n2127), .A4(n2126), .ZN(n2135)
         );
  OAI22_X1 U2271 ( .A1(n286), .A2(n2252), .B1(n574), .B2(n2265), .ZN(n2133) );
  OAI22_X1 U2272 ( .A1(n606), .A2(n2250), .B1(n254), .B2(n2263), .ZN(n2132) );
  OAI22_X1 U2273 ( .A1(n990), .A2(n2258), .B1(n766), .B2(n2276), .ZN(n2131) );
  OAI22_X1 U2274 ( .A1(n702), .A2(n2262), .B1(n414), .B2(n2270), .ZN(n2130) );
  NOR4_X1 U2275 ( .A1(n2133), .A2(n2132), .A3(n2131), .A4(n2130), .ZN(n2134)
         );
  NAND4_X1 U2276 ( .A1(n2137), .A2(n2136), .A3(n2135), .A4(n2134), .ZN(n2138)
         );
  AOI22_X1 U2277 ( .A1(n1680), .A2(n2138), .B1(n2281), .B2(lo_out[29]), .ZN(
        n2139) );
  OAI21_X1 U2278 ( .B1(n2283), .B2(n1646), .A(n2139), .ZN(rp1[29]) );
  NOR2_X1 U2279 ( .A1(n927), .A2(n2272), .ZN(n2143) );
  OAI22_X1 U2280 ( .A1(n575), .A2(n2265), .B1(n639), .B2(n2271), .ZN(n2142) );
  OAI22_X1 U2281 ( .A1(n671), .A2(n2278), .B1(n735), .B2(n2269), .ZN(n2141) );
  OAI22_X1 U2282 ( .A1(n511), .A2(n2259), .B1(n127), .B2(n2274), .ZN(n2140) );
  NOR4_X1 U2283 ( .A1(n2143), .A2(n2142), .A3(n2141), .A4(n2140), .ZN(n2159)
         );
  OAI22_X1 U2284 ( .A1(n191), .A2(n2257), .B1(n415), .B2(n2270), .ZN(n2147) );
  OAI22_X1 U2285 ( .A1(n351), .A2(n2256), .B1(n703), .B2(n2262), .ZN(n2146) );
  OAI22_X1 U2286 ( .A1(n447), .A2(n2267), .B1(n479), .B2(n2268), .ZN(n2145) );
  OAI22_X1 U2287 ( .A1(n831), .A2(n2273), .B1(n223), .B2(n2266), .ZN(n2144) );
  NOR4_X1 U2288 ( .A1(n2147), .A2(n2146), .A3(n2145), .A4(n2144), .ZN(n2158)
         );
  OAI22_X1 U2289 ( .A1(n799), .A2(n2279), .B1(n767), .B2(n2276), .ZN(n2151) );
  OAI22_X1 U2290 ( .A1(n543), .A2(n2253), .B1(n991), .B2(n2258), .ZN(n2150) );
  OAI22_X1 U2291 ( .A1(n959), .A2(n2277), .B1(n255), .B2(n2263), .ZN(n2149) );
  OAI22_X1 U2292 ( .A1(n383), .A2(n2260), .B1(n319), .B2(n2280), .ZN(n2148) );
  NOR4_X1 U2293 ( .A1(n2151), .A2(n2150), .A3(n2149), .A4(n2148), .ZN(n2157)
         );
  OAI22_X1 U2294 ( .A1(n31), .A2(n2264), .B1(n63), .B2(n2255), .ZN(n2155) );
  OAI22_X1 U2295 ( .A1(n895), .A2(n2275), .B1(n863), .B2(n2261), .ZN(n2154) );
  OAI22_X1 U2296 ( .A1(n287), .A2(n2252), .B1(n95), .B2(n2251), .ZN(n2153) );
  OAI22_X1 U2297 ( .A1(n159), .A2(n1677), .B1(n607), .B2(n2250), .ZN(n2152) );
  NOR4_X1 U2298 ( .A1(n2155), .A2(n2154), .A3(n2153), .A4(n2152), .ZN(n2156)
         );
  NAND4_X1 U2299 ( .A1(n2159), .A2(n2158), .A3(n2157), .A4(n2156), .ZN(n2160)
         );
  AOI22_X1 U2300 ( .A1(n1680), .A2(n2160), .B1(n2281), .B2(lo_out[30]), .ZN(
        n2161) );
  OAI21_X1 U2301 ( .B1(n2283), .B2(n1654), .A(n2161), .ZN(rp1[30]) );
  NOR2_X1 U2302 ( .A1(n192), .A2(n2257), .ZN(n2165) );
  OAI22_X1 U2303 ( .A1(n288), .A2(n2252), .B1(n352), .B2(n2256), .ZN(n2164) );
  OAI22_X1 U2304 ( .A1(n768), .A2(n2276), .B1(n96), .B2(n2251), .ZN(n2163) );
  OAI22_X1 U2305 ( .A1(n384), .A2(n2260), .B1(n256), .B2(n2263), .ZN(n2162) );
  NOR4_X1 U2306 ( .A1(n2165), .A2(n2164), .A3(n2163), .A4(n2162), .ZN(n2181)
         );
  OAI22_X1 U2307 ( .A1(n160), .A2(n1677), .B1(n928), .B2(n2272), .ZN(n2169) );
  OAI22_X1 U2308 ( .A1(n480), .A2(n2268), .B1(n128), .B2(n2274), .ZN(n2168) );
  OAI22_X1 U2309 ( .A1(n736), .A2(n2269), .B1(n32), .B2(n2264), .ZN(n2167) );
  OAI22_X1 U2310 ( .A1(n832), .A2(n2273), .B1(n448), .B2(n2267), .ZN(n2166) );
  NOR4_X1 U2311 ( .A1(n2169), .A2(n2168), .A3(n2167), .A4(n2166), .ZN(n2180)
         );
  OAI22_X1 U2312 ( .A1(n544), .A2(n2253), .B1(n416), .B2(n2270), .ZN(n2173) );
  OAI22_X1 U2313 ( .A1(n864), .A2(n2261), .B1(n704), .B2(n2262), .ZN(n2172) );
  OAI22_X1 U2314 ( .A1(n672), .A2(n2278), .B1(n64), .B2(n2255), .ZN(n2171) );
  OAI22_X1 U2315 ( .A1(n992), .A2(n2258), .B1(n608), .B2(n2250), .ZN(n2170) );
  NOR4_X1 U2316 ( .A1(n2173), .A2(n2172), .A3(n2171), .A4(n2170), .ZN(n2179)
         );
  OAI22_X1 U2317 ( .A1(n320), .A2(n2280), .B1(n800), .B2(n2279), .ZN(n2177) );
  OAI22_X1 U2318 ( .A1(n224), .A2(n2266), .B1(n512), .B2(n2259), .ZN(n2176) );
  OAI22_X1 U2319 ( .A1(n576), .A2(n2265), .B1(n896), .B2(n2275), .ZN(n2175) );
  OAI22_X1 U2320 ( .A1(n640), .A2(n1678), .B1(n960), .B2(n2277), .ZN(n2174) );
  NOR4_X1 U2321 ( .A1(n2177), .A2(n2176), .A3(n2175), .A4(n2174), .ZN(n2178)
         );
  NAND4_X1 U2322 ( .A1(n2181), .A2(n2180), .A3(n2179), .A4(n2178), .ZN(n2182)
         );
  AOI22_X1 U2323 ( .A1(n1680), .A2(n2182), .B1(n1679), .B2(lo_out[31]), .ZN(
        n2183) );
  OAI21_X1 U2324 ( .B1(n2283), .B2(n1647), .A(n2183), .ZN(rp1[31]) );
  NOR2_X1 U2325 ( .A1(n196), .A2(n2266), .ZN(n2187) );
  OAI22_X1 U2326 ( .A1(n708), .A2(n2269), .B1(n964), .B2(n2258), .ZN(n2186) );
  OAI22_X1 U2327 ( .A1(n292), .A2(n2280), .B1(n836), .B2(n2261), .ZN(n2185) );
  OAI22_X1 U2328 ( .A1(n868), .A2(n2275), .B1(n36), .B2(n2255), .ZN(n2184) );
  NOR4_X1 U2329 ( .A1(n2187), .A2(n2186), .A3(n2185), .A4(n2184), .ZN(n2203)
         );
  OAI22_X1 U2330 ( .A1(n164), .A2(n2257), .B1(n516), .B2(n2253), .ZN(n2191) );
  OAI22_X1 U2331 ( .A1(n740), .A2(n2276), .B1(n580), .B2(n2250), .ZN(n2190) );
  OAI22_X1 U2332 ( .A1(n324), .A2(n2256), .B1(n548), .B2(n2265), .ZN(n2189) );
  OAI22_X1 U2333 ( .A1(n772), .A2(n2279), .B1(n804), .B2(n2273), .ZN(n2188) );
  NOR4_X1 U2334 ( .A1(n2191), .A2(n2190), .A3(n2189), .A4(n2188), .ZN(n2202)
         );
  OAI22_X1 U2335 ( .A1(n932), .A2(n2277), .B1(n388), .B2(n2270), .ZN(n2195) );
  OAI22_X1 U2336 ( .A1(n4), .A2(n2264), .B1(n356), .B2(n2260), .ZN(n2194) );
  OAI22_X1 U2337 ( .A1(n900), .A2(n2272), .B1(n612), .B2(n1678), .ZN(n2193) );
  OAI22_X1 U2338 ( .A1(n228), .A2(n2263), .B1(n260), .B2(n2252), .ZN(n2192) );
  NOR4_X1 U2339 ( .A1(n2195), .A2(n2194), .A3(n2193), .A4(n2192), .ZN(n2201)
         );
  OAI22_X1 U2340 ( .A1(n452), .A2(n2268), .B1(n100), .B2(n2274), .ZN(n2199) );
  OAI22_X1 U2341 ( .A1(n484), .A2(n2259), .B1(n132), .B2(n2254), .ZN(n2198) );
  OAI22_X1 U2342 ( .A1(n420), .A2(n2267), .B1(n676), .B2(n2262), .ZN(n2197) );
  OAI22_X1 U2343 ( .A1(n644), .A2(n2278), .B1(n68), .B2(n2251), .ZN(n2196) );
  NOR4_X1 U2344 ( .A1(n2199), .A2(n2198), .A3(n2197), .A4(n2196), .ZN(n2200)
         );
  NAND4_X1 U2345 ( .A1(n2203), .A2(n2202), .A3(n2201), .A4(n2200), .ZN(n2204)
         );
  AOI22_X1 U2346 ( .A1(n1680), .A2(n2204), .B1(n1679), .B2(lo_out[3]), .ZN(
        n2205) );
  OAI21_X1 U2347 ( .B1(n2283), .B2(n1648), .A(n2205), .ZN(rp1[3]) );
  NOR2_X1 U2348 ( .A1(n581), .A2(n2250), .ZN(n2209) );
  OAI22_X1 U2349 ( .A1(n741), .A2(n2276), .B1(n101), .B2(n2274), .ZN(n2208) );
  OAI22_X1 U2350 ( .A1(n261), .A2(n2252), .B1(n389), .B2(n2270), .ZN(n2207) );
  OAI22_X1 U2351 ( .A1(n69), .A2(n2251), .B1(n645), .B2(n2278), .ZN(n2206) );
  NOR4_X1 U2352 ( .A1(n2209), .A2(n2208), .A3(n2207), .A4(n2206), .ZN(n2225)
         );
  OAI22_X1 U2353 ( .A1(n517), .A2(n2253), .B1(n805), .B2(n2273), .ZN(n2213) );
  OAI22_X1 U2354 ( .A1(n485), .A2(n2259), .B1(n293), .B2(n2280), .ZN(n2212) );
  OAI22_X1 U2355 ( .A1(n325), .A2(n2256), .B1(n869), .B2(n2275), .ZN(n2211) );
  OAI22_X1 U2356 ( .A1(n773), .A2(n2279), .B1(n197), .B2(n2266), .ZN(n2210) );
  NOR4_X1 U2357 ( .A1(n2213), .A2(n2212), .A3(n2211), .A4(n2210), .ZN(n2224)
         );
  OAI22_X1 U2358 ( .A1(n5), .A2(n2264), .B1(n837), .B2(n2261), .ZN(n2217) );
  OAI22_X1 U2359 ( .A1(n357), .A2(n2260), .B1(n677), .B2(n2262), .ZN(n2216) );
  OAI22_X1 U2360 ( .A1(n933), .A2(n2277), .B1(n709), .B2(n2269), .ZN(n2215) );
  OAI22_X1 U2361 ( .A1(n613), .A2(n1678), .B1(n133), .B2(n2254), .ZN(n2214) );
  NOR4_X1 U2362 ( .A1(n2217), .A2(n2216), .A3(n2215), .A4(n2214), .ZN(n2223)
         );
  OAI22_X1 U2363 ( .A1(n965), .A2(n2258), .B1(n37), .B2(n2255), .ZN(n2221) );
  OAI22_X1 U2364 ( .A1(n549), .A2(n2265), .B1(n421), .B2(n2267), .ZN(n2220) );
  OAI22_X1 U2365 ( .A1(n165), .A2(n2257), .B1(n453), .B2(n2268), .ZN(n2219) );
  OAI22_X1 U2366 ( .A1(n229), .A2(n2263), .B1(n901), .B2(n2272), .ZN(n2218) );
  NOR4_X1 U2367 ( .A1(n2221), .A2(n2220), .A3(n2219), .A4(n2218), .ZN(n2222)
         );
  NAND4_X1 U2368 ( .A1(n2225), .A2(n2224), .A3(n2223), .A4(n2222), .ZN(n2226)
         );
  AOI22_X1 U2369 ( .A1(n1680), .A2(n2226), .B1(n1679), .B2(lo_out[4]), .ZN(
        n2227) );
  OAI21_X1 U2370 ( .B1(n2283), .B2(n1649), .A(n2227), .ZN(rp1[4]) );
  NOR2_X1 U2371 ( .A1(n935), .A2(n2277), .ZN(n2231) );
  OAI22_X1 U2372 ( .A1(n135), .A2(n1677), .B1(n423), .B2(n2267), .ZN(n2230) );
  OAI22_X1 U2373 ( .A1(n7), .A2(n2264), .B1(n839), .B2(n2261), .ZN(n2229) );
  OAI22_X1 U2374 ( .A1(n903), .A2(n2272), .B1(n199), .B2(n2266), .ZN(n2228) );
  NOR4_X1 U2375 ( .A1(n2231), .A2(n2230), .A3(n2229), .A4(n2228), .ZN(n2247)
         );
  OAI22_X1 U2376 ( .A1(n327), .A2(n2256), .B1(n871), .B2(n2275), .ZN(n2235) );
  OAI22_X1 U2377 ( .A1(n615), .A2(n1678), .B1(n487), .B2(n2259), .ZN(n2234) );
  OAI22_X1 U2378 ( .A1(n231), .A2(n2263), .B1(n71), .B2(n2251), .ZN(n2233) );
  OAI22_X1 U2379 ( .A1(n391), .A2(n2270), .B1(n295), .B2(n2280), .ZN(n2232) );
  NOR4_X1 U2380 ( .A1(n2235), .A2(n2234), .A3(n2233), .A4(n2232), .ZN(n2246)
         );
  OAI22_X1 U2381 ( .A1(n647), .A2(n2278), .B1(n711), .B2(n2269), .ZN(n2239) );
  OAI22_X1 U2382 ( .A1(n39), .A2(n2255), .B1(n359), .B2(n2260), .ZN(n2238) );
  OAI22_X1 U2383 ( .A1(n167), .A2(n2257), .B1(n455), .B2(n2268), .ZN(n2237) );
  OAI22_X1 U2384 ( .A1(n807), .A2(n2273), .B1(n103), .B2(n2274), .ZN(n2236) );
  NOR4_X1 U2385 ( .A1(n2239), .A2(n2238), .A3(n2237), .A4(n2236), .ZN(n2245)
         );
  OAI22_X1 U2386 ( .A1(n263), .A2(n2252), .B1(n519), .B2(n2253), .ZN(n2243) );
  OAI22_X1 U2387 ( .A1(n551), .A2(n2265), .B1(n743), .B2(n2276), .ZN(n2242) );
  OAI22_X1 U2388 ( .A1(n775), .A2(n2279), .B1(n679), .B2(n2262), .ZN(n2241) );
  OAI22_X1 U2389 ( .A1(n967), .A2(n2258), .B1(n583), .B2(n2250), .ZN(n2240) );
  NOR4_X1 U2390 ( .A1(n2243), .A2(n2242), .A3(n2241), .A4(n2240), .ZN(n2244)
         );
  NAND4_X1 U2391 ( .A1(n2247), .A2(n2246), .A3(n2245), .A4(n2244), .ZN(n2248)
         );
  AOI22_X1 U2392 ( .A1(n1680), .A2(n2248), .B1(n1679), .B2(lo_out[6]), .ZN(
        n2249) );
  OAI21_X1 U2393 ( .B1(n2283), .B2(n1624), .A(n2249), .ZN(rp1[6]) );
  NOR2_X1 U2394 ( .A1(rp2_out_sel[1]), .A2(n2284), .ZN(n3786) );
  NOR2_X1 U2395 ( .A1(rp2_out_sel[1]), .A2(rp2_out_sel[0]), .ZN(n3785) );
  AND2_X1 U2396 ( .A1(rp2_addr[1]), .A2(rp2_addr[2]), .ZN(n2307) );
  INV_X1 U2397 ( .A(rp2_addr[3]), .ZN(n2285) );
  NOR3_X1 U2398 ( .A1(rp2_addr[0]), .A2(rp2_addr[4]), .A3(n2285), .ZN(n2298)
         );
  NOR2_X1 U2399 ( .A1(n417), .A2(n3760), .ZN(n2291) );
  INV_X1 U2400 ( .A(rp2_addr[0]), .ZN(n2293) );
  NOR3_X1 U2401 ( .A1(rp2_addr[3]), .A2(rp2_addr[4]), .A3(n2293), .ZN(n2304)
         );
  NOR2_X1 U2402 ( .A1(rp2_addr[1]), .A2(rp2_addr[2]), .ZN(n2311) );
  NAND2_X1 U2403 ( .A1(rp2_addr[3]), .A2(rp2_addr[4]), .ZN(n2292) );
  NOR2_X1 U2404 ( .A1(rp2_addr[0]), .A2(n2292), .ZN(n2305) );
  OAI22_X1 U2405 ( .A1(n193), .A2(n3758), .B1(n737), .B2(n3768), .ZN(n2290) );
  INV_X1 U2406 ( .A(rp2_addr[2]), .ZN(n2287) );
  NOR2_X1 U2407 ( .A1(rp2_addr[1]), .A2(n2287), .ZN(n2310) );
  NOR3_X1 U2408 ( .A1(rp2_addr[4]), .A2(n2285), .A3(n2293), .ZN(n2313) );
  NAND2_X1 U2409 ( .A1(n2310), .A2(n2313), .ZN(n3780) );
  INV_X1 U2410 ( .A(rp2_addr[4]), .ZN(n2286) );
  NOR3_X1 U2411 ( .A1(rp2_addr[3]), .A2(n2293), .A3(n2286), .ZN(n2299) );
  OAI22_X1 U2412 ( .A1(n385), .A2(n3780), .B1(n705), .B2(n3762), .ZN(n2289) );
  NAND2_X1 U2413 ( .A1(n2304), .A2(n2310), .ZN(n3769) );
  NOR3_X1 U2414 ( .A1(rp2_addr[0]), .A2(rp2_addr[3]), .A3(n2286), .ZN(n2306)
         );
  AND2_X1 U2415 ( .A1(n2287), .A2(rp2_addr[1]), .ZN(n2312) );
  OAI22_X1 U2416 ( .A1(n129), .A2(n1682), .B1(n545), .B2(n3782), .ZN(n2288) );
  NOR4_X1 U2417 ( .A1(n2291), .A2(n2290), .A3(n2289), .A4(n2288), .ZN(n2321)
         );
  NOR2_X1 U2418 ( .A1(n2293), .A2(n2292), .ZN(n2308) );
  OAI22_X1 U2419 ( .A1(n833), .A2(n3767), .B1(n929), .B2(n3784), .ZN(n2297) );
  NAND2_X1 U2420 ( .A1(n2310), .A2(n2306), .ZN(n3755) );
  OAI22_X1 U2421 ( .A1(n641), .A2(n3756), .B1(n609), .B2(n3755), .ZN(n2296) );
  OAI22_X1 U2422 ( .A1(n577), .A2(n3759), .B1(n353), .B2(n3776), .ZN(n2295) );
  OAI22_X1 U2423 ( .A1(n225), .A2(n3781), .B1(n481), .B2(n3757), .ZN(n2294) );
  NOR4_X1 U2424 ( .A1(n2297), .A2(n2296), .A3(n2295), .A4(n2294), .ZN(n2320)
         );
  NOR3_X1 U2425 ( .A1(rp2_addr[0]), .A2(rp2_addr[3]), .A3(rp2_addr[4]), .ZN(
        n2309) );
  OAI22_X1 U2426 ( .A1(n33), .A2(n3773), .B1(n961), .B2(n3771), .ZN(n2303) );
  OAI22_X1 U2427 ( .A1(n1), .A2(n3770), .B1(n801), .B2(n3754), .ZN(n2302) );
  OAI22_X1 U2428 ( .A1(n289), .A2(n3764), .B1(n449), .B2(n3766), .ZN(n2301) );
  OAI22_X1 U2429 ( .A1(n513), .A2(n3779), .B1(n897), .B2(n3783), .ZN(n2300) );
  NOR4_X1 U2430 ( .A1(n2303), .A2(n2302), .A3(n2301), .A4(n2300), .ZN(n2319)
         );
  OAI22_X1 U2431 ( .A1(n65), .A2(n3763), .B1(n865), .B2(n3778), .ZN(n2317) );
  OAI22_X1 U2432 ( .A1(n161), .A2(n3761), .B1(n673), .B2(n3765), .ZN(n2316) );
  OAI22_X1 U2433 ( .A1(n769), .A2(n3772), .B1(n97), .B2(n3774), .ZN(n2315) );
  OAI22_X1 U2434 ( .A1(n257), .A2(n3775), .B1(n321), .B2(n3777), .ZN(n2314) );
  NOR4_X1 U2435 ( .A1(n2317), .A2(n2316), .A3(n2315), .A4(n2314), .ZN(n2318)
         );
  NAND4_X1 U2436 ( .A1(n2321), .A2(n2320), .A3(n2319), .A4(n2318), .ZN(n2322)
         );
  AOI22_X1 U2437 ( .A1(lo_out[0]), .A2(n1685), .B1(n3785), .B2(n2322), .ZN(
        n2323) );
  OAI21_X1 U2438 ( .B1(n1628), .B2(n3787), .A(n2323), .ZN(rp2[0]) );
  NOR2_X1 U2439 ( .A1(n209), .A2(n3758), .ZN(n2327) );
  OAI22_X1 U2440 ( .A1(n369), .A2(n3776), .B1(n465), .B2(n3766), .ZN(n2326) );
  OAI22_X1 U2441 ( .A1(n753), .A2(n3768), .B1(n593), .B2(n3759), .ZN(n2325) );
  OAI22_X1 U2442 ( .A1(n433), .A2(n3760), .B1(n177), .B2(n3761), .ZN(n2324) );
  NOR4_X1 U2443 ( .A1(n2327), .A2(n2326), .A3(n2325), .A4(n2324), .ZN(n2343)
         );
  OAI22_X1 U2444 ( .A1(n721), .A2(n3762), .B1(n785), .B2(n3772), .ZN(n2331) );
  OAI22_X1 U2445 ( .A1(n849), .A2(n3767), .B1(n49), .B2(n3773), .ZN(n2330) );
  OAI22_X1 U2446 ( .A1(n561), .A2(n3782), .B1(n689), .B2(n3765), .ZN(n2329) );
  OAI22_X1 U2447 ( .A1(n81), .A2(n3763), .B1(n657), .B2(n3756), .ZN(n2328) );
  NOR4_X1 U2448 ( .A1(n2331), .A2(n2330), .A3(n2329), .A4(n2328), .ZN(n2342)
         );
  OAI22_X1 U2449 ( .A1(n945), .A2(n3784), .B1(n817), .B2(n3754), .ZN(n2335) );
  OAI22_X1 U2450 ( .A1(n977), .A2(n3771), .B1(n401), .B2(n1683), .ZN(n2334) );
  OAI22_X1 U2451 ( .A1(n17), .A2(n3770), .B1(n913), .B2(n3783), .ZN(n2333) );
  OAI22_X1 U2452 ( .A1(n337), .A2(n3777), .B1(n625), .B2(n1681), .ZN(n2332) );
  NOR4_X1 U2453 ( .A1(n2335), .A2(n2334), .A3(n2333), .A4(n2332), .ZN(n2341)
         );
  OAI22_X1 U2454 ( .A1(n113), .A2(n3774), .B1(n145), .B2(n3769), .ZN(n2339) );
  OAI22_X1 U2455 ( .A1(n881), .A2(n3778), .B1(n273), .B2(n3775), .ZN(n2338) );
  OAI22_X1 U2456 ( .A1(n529), .A2(n3779), .B1(n305), .B2(n3764), .ZN(n2337) );
  OAI22_X1 U2457 ( .A1(n497), .A2(n3757), .B1(n241), .B2(n3781), .ZN(n2336) );
  NOR4_X1 U2458 ( .A1(n2339), .A2(n2338), .A3(n2337), .A4(n2336), .ZN(n2340)
         );
  NAND4_X1 U2459 ( .A1(n2343), .A2(n2342), .A3(n2341), .A4(n2340), .ZN(n2344)
         );
  AOI22_X1 U2460 ( .A1(lo_out[16]), .A2(n1685), .B1(n1684), .B2(n2344), .ZN(
        n2345) );
  OAI21_X1 U2461 ( .B1(n1635), .B2(n3787), .A(n2345), .ZN(rp2[16]) );
  NOR2_X1 U2462 ( .A1(n434), .A2(n3760), .ZN(n2349) );
  OAI22_X1 U2463 ( .A1(n530), .A2(n3779), .B1(n306), .B2(n3764), .ZN(n2348) );
  OAI22_X1 U2464 ( .A1(n82), .A2(n3763), .B1(n658), .B2(n3756), .ZN(n2347) );
  OAI22_X1 U2465 ( .A1(n754), .A2(n3768), .B1(n786), .B2(n3772), .ZN(n2346) );
  NOR4_X1 U2466 ( .A1(n2349), .A2(n2348), .A3(n2347), .A4(n2346), .ZN(n2365)
         );
  OAI22_X1 U2467 ( .A1(n370), .A2(n3776), .B1(n466), .B2(n3766), .ZN(n2353) );
  OAI22_X1 U2468 ( .A1(n50), .A2(n3773), .B1(n338), .B2(n3777), .ZN(n2352) );
  OAI22_X1 U2469 ( .A1(n818), .A2(n3754), .B1(n242), .B2(n3781), .ZN(n2351) );
  OAI22_X1 U2470 ( .A1(n626), .A2(n3755), .B1(n498), .B2(n3757), .ZN(n2350) );
  NOR4_X1 U2471 ( .A1(n2353), .A2(n2352), .A3(n2351), .A4(n2350), .ZN(n2364)
         );
  OAI22_X1 U2472 ( .A1(n402), .A2(n1683), .B1(n178), .B2(n3761), .ZN(n2357) );
  OAI22_X1 U2473 ( .A1(n946), .A2(n3784), .B1(n18), .B2(n3770), .ZN(n2356) );
  OAI22_X1 U2474 ( .A1(n978), .A2(n3771), .B1(n882), .B2(n3778), .ZN(n2355) );
  OAI22_X1 U2475 ( .A1(n210), .A2(n3758), .B1(n562), .B2(n3782), .ZN(n2354) );
  NOR4_X1 U2476 ( .A1(n2357), .A2(n2356), .A3(n2355), .A4(n2354), .ZN(n2363)
         );
  OAI22_X1 U2477 ( .A1(n850), .A2(n3767), .B1(n722), .B2(n3762), .ZN(n2361) );
  OAI22_X1 U2478 ( .A1(n690), .A2(n3765), .B1(n914), .B2(n3783), .ZN(n2360) );
  OAI22_X1 U2479 ( .A1(n146), .A2(n1682), .B1(n274), .B2(n3775), .ZN(n2359) );
  OAI22_X1 U2480 ( .A1(n114), .A2(n3774), .B1(n594), .B2(n3759), .ZN(n2358) );
  NOR4_X1 U2481 ( .A1(n2361), .A2(n2360), .A3(n2359), .A4(n2358), .ZN(n2362)
         );
  NAND4_X1 U2482 ( .A1(n2365), .A2(n2364), .A3(n2363), .A4(n2362), .ZN(n2366)
         );
  AOI22_X1 U2483 ( .A1(lo_out[17]), .A2(n1685), .B1(n3785), .B2(n2366), .ZN(
        n2367) );
  OAI21_X1 U2484 ( .B1(n1650), .B2(n3787), .A(n2367), .ZN(rp2[17]) );
  NOR2_X1 U2485 ( .A1(n275), .A2(n3775), .ZN(n2371) );
  OAI22_X1 U2486 ( .A1(n851), .A2(n3767), .B1(n307), .B2(n3764), .ZN(n2370) );
  OAI22_X1 U2487 ( .A1(n691), .A2(n3765), .B1(n403), .B2(n1683), .ZN(n2369) );
  OAI22_X1 U2488 ( .A1(n659), .A2(n3756), .B1(n371), .B2(n3776), .ZN(n2368) );
  NOR4_X1 U2489 ( .A1(n2371), .A2(n2370), .A3(n2369), .A4(n2368), .ZN(n2387)
         );
  OAI22_X1 U2490 ( .A1(n915), .A2(n3783), .B1(n787), .B2(n3772), .ZN(n2375) );
  OAI22_X1 U2491 ( .A1(n595), .A2(n3759), .B1(n467), .B2(n3766), .ZN(n2374) );
  OAI22_X1 U2492 ( .A1(n339), .A2(n3777), .B1(n947), .B2(n3784), .ZN(n2373) );
  OAI22_X1 U2493 ( .A1(n115), .A2(n3774), .B1(n147), .B2(n3769), .ZN(n2372) );
  NOR4_X1 U2494 ( .A1(n2375), .A2(n2374), .A3(n2373), .A4(n2372), .ZN(n2386)
         );
  OAI22_X1 U2495 ( .A1(n979), .A2(n3771), .B1(n499), .B2(n3757), .ZN(n2379) );
  OAI22_X1 U2496 ( .A1(n563), .A2(n3782), .B1(n627), .B2(n1681), .ZN(n2378) );
  OAI22_X1 U2497 ( .A1(n243), .A2(n3781), .B1(n211), .B2(n3758), .ZN(n2377) );
  OAI22_X1 U2498 ( .A1(n531), .A2(n3779), .B1(n19), .B2(n3770), .ZN(n2376) );
  NOR4_X1 U2499 ( .A1(n2379), .A2(n2378), .A3(n2377), .A4(n2376), .ZN(n2385)
         );
  OAI22_X1 U2500 ( .A1(n179), .A2(n3761), .B1(n819), .B2(n3754), .ZN(n2383) );
  OAI22_X1 U2501 ( .A1(n723), .A2(n3762), .B1(n755), .B2(n3768), .ZN(n2382) );
  OAI22_X1 U2502 ( .A1(n883), .A2(n3778), .B1(n51), .B2(n3773), .ZN(n2381) );
  OAI22_X1 U2503 ( .A1(n83), .A2(n3763), .B1(n435), .B2(n3760), .ZN(n2380) );
  NOR4_X1 U2504 ( .A1(n2383), .A2(n2382), .A3(n2381), .A4(n2380), .ZN(n2384)
         );
  NAND4_X1 U2505 ( .A1(n2387), .A2(n2386), .A3(n2385), .A4(n2384), .ZN(n2388)
         );
  AOI22_X1 U2506 ( .A1(lo_out[18]), .A2(n1685), .B1(n1684), .B2(n2388), .ZN(
        n2389) );
  OAI21_X1 U2507 ( .B1(n1636), .B2(n3787), .A(n2389), .ZN(rp2[18]) );
  NOR2_X1 U2508 ( .A1(n564), .A2(n3782), .ZN(n2393) );
  OAI22_X1 U2509 ( .A1(n916), .A2(n3783), .B1(n84), .B2(n3763), .ZN(n2392) );
  OAI22_X1 U2510 ( .A1(n20), .A2(n3770), .B1(n724), .B2(n3762), .ZN(n2391) );
  OAI22_X1 U2511 ( .A1(n852), .A2(n3767), .B1(n52), .B2(n3773), .ZN(n2390) );
  NOR4_X1 U2512 ( .A1(n2393), .A2(n2392), .A3(n2391), .A4(n2390), .ZN(n2409)
         );
  OAI22_X1 U2513 ( .A1(n756), .A2(n3768), .B1(n500), .B2(n3757), .ZN(n2397) );
  OAI22_X1 U2514 ( .A1(n980), .A2(n3771), .B1(n820), .B2(n3754), .ZN(n2396) );
  OAI22_X1 U2515 ( .A1(n948), .A2(n3784), .B1(n340), .B2(n3777), .ZN(n2395) );
  OAI22_X1 U2516 ( .A1(n596), .A2(n3759), .B1(n468), .B2(n3766), .ZN(n2394) );
  NOR4_X1 U2517 ( .A1(n2397), .A2(n2396), .A3(n2395), .A4(n2394), .ZN(n2408)
         );
  OAI22_X1 U2518 ( .A1(n148), .A2(n3769), .B1(n212), .B2(n3758), .ZN(n2401) );
  OAI22_X1 U2519 ( .A1(n884), .A2(n3778), .B1(n244), .B2(n3781), .ZN(n2400) );
  OAI22_X1 U2520 ( .A1(n372), .A2(n3776), .B1(n180), .B2(n3761), .ZN(n2399) );
  OAI22_X1 U2521 ( .A1(n276), .A2(n3775), .B1(n116), .B2(n3774), .ZN(n2398) );
  NOR4_X1 U2522 ( .A1(n2401), .A2(n2400), .A3(n2399), .A4(n2398), .ZN(n2407)
         );
  OAI22_X1 U2523 ( .A1(n532), .A2(n3779), .B1(n660), .B2(n3756), .ZN(n2405) );
  OAI22_X1 U2524 ( .A1(n788), .A2(n3772), .B1(n436), .B2(n3760), .ZN(n2404) );
  OAI22_X1 U2525 ( .A1(n692), .A2(n3765), .B1(n404), .B2(n1683), .ZN(n2403) );
  OAI22_X1 U2526 ( .A1(n628), .A2(n1681), .B1(n308), .B2(n3764), .ZN(n2402) );
  NOR4_X1 U2527 ( .A1(n2405), .A2(n2404), .A3(n2403), .A4(n2402), .ZN(n2406)
         );
  NAND4_X1 U2528 ( .A1(n2409), .A2(n2408), .A3(n2407), .A4(n2406), .ZN(n2410)
         );
  AOI22_X1 U2529 ( .A1(lo_out[19]), .A2(n1685), .B1(n1684), .B2(n2410), .ZN(
        n2411) );
  OAI21_X1 U2530 ( .B1(n1637), .B2(n3787), .A(n2411), .ZN(rp2[19]) );
  NOR2_X1 U2531 ( .A1(n386), .A2(n1683), .ZN(n2415) );
  OAI22_X1 U2532 ( .A1(n802), .A2(n3754), .B1(n674), .B2(n3765), .ZN(n2414) );
  OAI22_X1 U2533 ( .A1(n706), .A2(n3762), .B1(n226), .B2(n3781), .ZN(n2413) );
  OAI22_X1 U2534 ( .A1(n290), .A2(n3764), .B1(n258), .B2(n3775), .ZN(n2412) );
  NOR4_X1 U2535 ( .A1(n2415), .A2(n2414), .A3(n2413), .A4(n2412), .ZN(n2431)
         );
  OAI22_X1 U2536 ( .A1(n962), .A2(n3771), .B1(n162), .B2(n3761), .ZN(n2419) );
  OAI22_X1 U2537 ( .A1(n34), .A2(n3773), .B1(n642), .B2(n3756), .ZN(n2418) );
  OAI22_X1 U2538 ( .A1(n130), .A2(n3769), .B1(n578), .B2(n3759), .ZN(n2417) );
  OAI22_X1 U2539 ( .A1(n66), .A2(n3763), .B1(n898), .B2(n3783), .ZN(n2416) );
  NOR4_X1 U2540 ( .A1(n2419), .A2(n2418), .A3(n2417), .A4(n2416), .ZN(n2430)
         );
  OAI22_X1 U2541 ( .A1(n834), .A2(n3767), .B1(n194), .B2(n3758), .ZN(n2423) );
  OAI22_X1 U2542 ( .A1(n354), .A2(n3776), .B1(n98), .B2(n3774), .ZN(n2422) );
  OAI22_X1 U2543 ( .A1(n514), .A2(n3779), .B1(n450), .B2(n3766), .ZN(n2421) );
  OAI22_X1 U2544 ( .A1(n2), .A2(n3770), .B1(n930), .B2(n3784), .ZN(n2420) );
  NOR4_X1 U2545 ( .A1(n2423), .A2(n2422), .A3(n2421), .A4(n2420), .ZN(n2429)
         );
  OAI22_X1 U2546 ( .A1(n770), .A2(n3772), .B1(n610), .B2(n1681), .ZN(n2427) );
  OAI22_X1 U2547 ( .A1(n546), .A2(n3782), .B1(n738), .B2(n3768), .ZN(n2426) );
  OAI22_X1 U2548 ( .A1(n482), .A2(n3757), .B1(n322), .B2(n3777), .ZN(n2425) );
  OAI22_X1 U2549 ( .A1(n866), .A2(n3778), .B1(n418), .B2(n3760), .ZN(n2424) );
  NOR4_X1 U2550 ( .A1(n2427), .A2(n2426), .A3(n2425), .A4(n2424), .ZN(n2428)
         );
  NAND4_X1 U2551 ( .A1(n2431), .A2(n2430), .A3(n2429), .A4(n2428), .ZN(n2432)
         );
  AOI22_X1 U2552 ( .A1(lo_out[1]), .A2(n1685), .B1(n3785), .B2(n2432), .ZN(
        n2433) );
  OAI21_X1 U2553 ( .B1(n1651), .B2(n3787), .A(n2433), .ZN(rp2[1]) );
  NOR2_X1 U2554 ( .A1(n405), .A2(n1683), .ZN(n2437) );
  OAI22_X1 U2555 ( .A1(n373), .A2(n3776), .B1(n437), .B2(n3760), .ZN(n2436) );
  OAI22_X1 U2556 ( .A1(n981), .A2(n3771), .B1(n309), .B2(n3764), .ZN(n2435) );
  OAI22_X1 U2557 ( .A1(n821), .A2(n3754), .B1(n725), .B2(n3762), .ZN(n2434) );
  NOR4_X1 U2558 ( .A1(n2437), .A2(n2436), .A3(n2435), .A4(n2434), .ZN(n2453)
         );
  OAI22_X1 U2559 ( .A1(n213), .A2(n3758), .B1(n85), .B2(n3763), .ZN(n2441) );
  OAI22_X1 U2560 ( .A1(n277), .A2(n3775), .B1(n501), .B2(n3757), .ZN(n2440) );
  OAI22_X1 U2561 ( .A1(n597), .A2(n3759), .B1(n629), .B2(n1681), .ZN(n2439) );
  OAI22_X1 U2562 ( .A1(n693), .A2(n3765), .B1(n533), .B2(n3779), .ZN(n2438) );
  NOR4_X1 U2563 ( .A1(n2441), .A2(n2440), .A3(n2439), .A4(n2438), .ZN(n2452)
         );
  OAI22_X1 U2564 ( .A1(n885), .A2(n3778), .B1(n757), .B2(n3768), .ZN(n2445) );
  OAI22_X1 U2565 ( .A1(n853), .A2(n3767), .B1(n53), .B2(n3773), .ZN(n2444) );
  OAI22_X1 U2566 ( .A1(n245), .A2(n3781), .B1(n789), .B2(n3772), .ZN(n2443) );
  OAI22_X1 U2567 ( .A1(n181), .A2(n3761), .B1(n469), .B2(n3766), .ZN(n2442) );
  NOR4_X1 U2568 ( .A1(n2445), .A2(n2444), .A3(n2443), .A4(n2442), .ZN(n2451)
         );
  OAI22_X1 U2569 ( .A1(n949), .A2(n3784), .B1(n661), .B2(n3756), .ZN(n2449) );
  OAI22_X1 U2570 ( .A1(n565), .A2(n3782), .B1(n117), .B2(n3774), .ZN(n2448) );
  OAI22_X1 U2571 ( .A1(n149), .A2(n3769), .B1(n341), .B2(n3777), .ZN(n2447) );
  OAI22_X1 U2572 ( .A1(n917), .A2(n3783), .B1(n21), .B2(n3770), .ZN(n2446) );
  NOR4_X1 U2573 ( .A1(n2449), .A2(n2448), .A3(n2447), .A4(n2446), .ZN(n2450)
         );
  NAND4_X1 U2574 ( .A1(n2453), .A2(n2452), .A3(n2451), .A4(n2450), .ZN(n2454)
         );
  AOI22_X1 U2575 ( .A1(lo_out[20]), .A2(n3786), .B1(n1684), .B2(n2454), .ZN(
        n2455) );
  OAI21_X1 U2576 ( .B1(n1638), .B2(n3787), .A(n2455), .ZN(rp2[20]) );
  NOR2_X1 U2577 ( .A1(n566), .A2(n3782), .ZN(n2459) );
  OAI22_X1 U2578 ( .A1(n598), .A2(n3759), .B1(n438), .B2(n3760), .ZN(n2458) );
  OAI22_X1 U2579 ( .A1(n822), .A2(n3754), .B1(n534), .B2(n3779), .ZN(n2457) );
  OAI22_X1 U2580 ( .A1(n470), .A2(n3766), .B1(n502), .B2(n3757), .ZN(n2456) );
  NOR4_X1 U2581 ( .A1(n2459), .A2(n2458), .A3(n2457), .A4(n2456), .ZN(n2475)
         );
  OAI22_X1 U2582 ( .A1(n278), .A2(n3775), .B1(n726), .B2(n3762), .ZN(n2463) );
  OAI22_X1 U2583 ( .A1(n86), .A2(n3763), .B1(n118), .B2(n3774), .ZN(n2462) );
  OAI22_X1 U2584 ( .A1(n950), .A2(n3784), .B1(n854), .B2(n3767), .ZN(n2461) );
  OAI22_X1 U2585 ( .A1(n758), .A2(n3768), .B1(n246), .B2(n3781), .ZN(n2460) );
  NOR4_X1 U2586 ( .A1(n2463), .A2(n2462), .A3(n2461), .A4(n2460), .ZN(n2474)
         );
  OAI22_X1 U2587 ( .A1(n918), .A2(n3783), .B1(n182), .B2(n3761), .ZN(n2467) );
  OAI22_X1 U2588 ( .A1(n214), .A2(n3758), .B1(n694), .B2(n3765), .ZN(n2466) );
  OAI22_X1 U2589 ( .A1(n630), .A2(n1681), .B1(n342), .B2(n3777), .ZN(n2465) );
  OAI22_X1 U2590 ( .A1(n310), .A2(n3764), .B1(n406), .B2(n1683), .ZN(n2464) );
  NOR4_X1 U2591 ( .A1(n2467), .A2(n2466), .A3(n2465), .A4(n2464), .ZN(n2473)
         );
  OAI22_X1 U2592 ( .A1(n886), .A2(n3778), .B1(n982), .B2(n3771), .ZN(n2471) );
  OAI22_X1 U2593 ( .A1(n662), .A2(n3756), .B1(n54), .B2(n3773), .ZN(n2470) );
  OAI22_X1 U2594 ( .A1(n22), .A2(n3770), .B1(n790), .B2(n3772), .ZN(n2469) );
  OAI22_X1 U2595 ( .A1(n374), .A2(n3776), .B1(n150), .B2(n1682), .ZN(n2468) );
  NOR4_X1 U2596 ( .A1(n2471), .A2(n2470), .A3(n2469), .A4(n2468), .ZN(n2472)
         );
  NAND4_X1 U2597 ( .A1(n2475), .A2(n2474), .A3(n2473), .A4(n2472), .ZN(n2476)
         );
  AOI22_X1 U2598 ( .A1(lo_out[21]), .A2(n3786), .B1(n1684), .B2(n2476), .ZN(
        n2477) );
  OAI21_X1 U2599 ( .B1(n1639), .B2(n3787), .A(n2477), .ZN(rp2[21]) );
  NOR2_X1 U2600 ( .A1(n951), .A2(n3784), .ZN(n2481) );
  OAI22_X1 U2601 ( .A1(n983), .A2(n3771), .B1(n343), .B2(n3777), .ZN(n2480) );
  OAI22_X1 U2602 ( .A1(n55), .A2(n3773), .B1(n919), .B2(n3783), .ZN(n2479) );
  OAI22_X1 U2603 ( .A1(n23), .A2(n3770), .B1(n311), .B2(n3764), .ZN(n2478) );
  NOR4_X1 U2604 ( .A1(n2481), .A2(n2480), .A3(n2479), .A4(n2478), .ZN(n2561)
         );
  OAI22_X1 U2605 ( .A1(n247), .A2(n3781), .B1(n823), .B2(n3754), .ZN(n2549) );
  OAI22_X1 U2606 ( .A1(n727), .A2(n3762), .B1(n599), .B2(n3759), .ZN(n2548) );
  OAI22_X1 U2607 ( .A1(n407), .A2(n3780), .B1(n471), .B2(n3766), .ZN(n2484) );
  OAI22_X1 U2608 ( .A1(n631), .A2(n1681), .B1(n439), .B2(n3760), .ZN(n2483) );
  NOR4_X1 U2609 ( .A1(n2549), .A2(n2548), .A3(n2484), .A4(n2483), .ZN(n2560)
         );
  OAI22_X1 U2610 ( .A1(n375), .A2(n3776), .B1(n279), .B2(n3775), .ZN(n2553) );
  OAI22_X1 U2611 ( .A1(n567), .A2(n3782), .B1(n535), .B2(n3779), .ZN(n2552) );
  OAI22_X1 U2612 ( .A1(n151), .A2(n3769), .B1(n791), .B2(n3772), .ZN(n2551) );
  OAI22_X1 U2613 ( .A1(n887), .A2(n3778), .B1(n503), .B2(n3757), .ZN(n2550) );
  NOR4_X1 U2614 ( .A1(n2553), .A2(n2552), .A3(n2551), .A4(n2550), .ZN(n2559)
         );
  OAI22_X1 U2615 ( .A1(n183), .A2(n3761), .B1(n119), .B2(n3774), .ZN(n2557) );
  OAI22_X1 U2616 ( .A1(n759), .A2(n3768), .B1(n87), .B2(n3763), .ZN(n2556) );
  OAI22_X1 U2617 ( .A1(n663), .A2(n3756), .B1(n695), .B2(n3765), .ZN(n2555) );
  OAI22_X1 U2618 ( .A1(n855), .A2(n3767), .B1(n215), .B2(n3758), .ZN(n2554) );
  NOR4_X1 U2619 ( .A1(n2557), .A2(n2556), .A3(n2555), .A4(n2554), .ZN(n2558)
         );
  NAND4_X1 U2620 ( .A1(n2561), .A2(n2560), .A3(n2559), .A4(n2558), .ZN(n2562)
         );
  AOI22_X1 U2621 ( .A1(lo_out[22]), .A2(n1685), .B1(n1684), .B2(n2562), .ZN(
        n2563) );
  OAI21_X1 U2622 ( .B1(n1640), .B2(n3787), .A(n2563), .ZN(rp2[22]) );
  NOR2_X1 U2623 ( .A1(n280), .A2(n3775), .ZN(n2567) );
  OAI22_X1 U2624 ( .A1(n632), .A2(n3755), .B1(n792), .B2(n3772), .ZN(n2566) );
  OAI22_X1 U2625 ( .A1(n216), .A2(n3758), .B1(n664), .B2(n3756), .ZN(n2565) );
  OAI22_X1 U2626 ( .A1(n120), .A2(n3774), .B1(n536), .B2(n3779), .ZN(n2564) );
  NOR4_X1 U2627 ( .A1(n2567), .A2(n2566), .A3(n2565), .A4(n2564), .ZN(n2583)
         );
  OAI22_X1 U2628 ( .A1(n728), .A2(n3762), .B1(n568), .B2(n3782), .ZN(n2571) );
  OAI22_X1 U2629 ( .A1(n920), .A2(n3783), .B1(n600), .B2(n3759), .ZN(n2570) );
  OAI22_X1 U2630 ( .A1(n952), .A2(n3784), .B1(n152), .B2(n1682), .ZN(n2569) );
  OAI22_X1 U2631 ( .A1(n56), .A2(n3773), .B1(n504), .B2(n3757), .ZN(n2568) );
  NOR4_X1 U2632 ( .A1(n2571), .A2(n2570), .A3(n2569), .A4(n2568), .ZN(n2582)
         );
  OAI22_X1 U2633 ( .A1(n344), .A2(n3777), .B1(n472), .B2(n3766), .ZN(n2575) );
  OAI22_X1 U2634 ( .A1(n440), .A2(n3760), .B1(n184), .B2(n3761), .ZN(n2574) );
  OAI22_X1 U2635 ( .A1(n856), .A2(n3767), .B1(n984), .B2(n3771), .ZN(n2573) );
  OAI22_X1 U2636 ( .A1(n24), .A2(n3770), .B1(n248), .B2(n3781), .ZN(n2572) );
  NOR4_X1 U2637 ( .A1(n2575), .A2(n2574), .A3(n2573), .A4(n2572), .ZN(n2581)
         );
  OAI22_X1 U2638 ( .A1(n824), .A2(n3754), .B1(n408), .B2(n3780), .ZN(n2579) );
  OAI22_X1 U2639 ( .A1(n312), .A2(n3764), .B1(n888), .B2(n3778), .ZN(n2578) );
  OAI22_X1 U2640 ( .A1(n760), .A2(n3768), .B1(n696), .B2(n3765), .ZN(n2577) );
  OAI22_X1 U2641 ( .A1(n376), .A2(n3776), .B1(n88), .B2(n3763), .ZN(n2576) );
  NOR4_X1 U2642 ( .A1(n2579), .A2(n2578), .A3(n2577), .A4(n2576), .ZN(n2580)
         );
  NAND4_X1 U2643 ( .A1(n2583), .A2(n2582), .A3(n2581), .A4(n2580), .ZN(n2584)
         );
  AOI22_X1 U2644 ( .A1(lo_out[23]), .A2(n1685), .B1(n3785), .B2(n2584), .ZN(
        n2585) );
  OAI21_X1 U2645 ( .B1(n1641), .B2(n3787), .A(n2585), .ZN(rp2[23]) );
  NOR2_X1 U2646 ( .A1(n889), .A2(n3778), .ZN(n2589) );
  OAI22_X1 U2647 ( .A1(n57), .A2(n3773), .B1(n185), .B2(n3761), .ZN(n2588) );
  OAI22_X1 U2648 ( .A1(n25), .A2(n3770), .B1(n409), .B2(n1683), .ZN(n2587) );
  OAI22_X1 U2649 ( .A1(n217), .A2(n3758), .B1(n953), .B2(n3784), .ZN(n2586) );
  NOR4_X1 U2650 ( .A1(n2589), .A2(n2588), .A3(n2587), .A4(n2586), .ZN(n2605)
         );
  OAI22_X1 U2651 ( .A1(n761), .A2(n3768), .B1(n985), .B2(n3771), .ZN(n2593) );
  OAI22_X1 U2652 ( .A1(n473), .A2(n3766), .B1(n441), .B2(n3760), .ZN(n2592) );
  OAI22_X1 U2653 ( .A1(n89), .A2(n3763), .B1(n153), .B2(n3769), .ZN(n2591) );
  OAI22_X1 U2654 ( .A1(n281), .A2(n3775), .B1(n825), .B2(n3754), .ZN(n2590) );
  NOR4_X1 U2655 ( .A1(n2593), .A2(n2592), .A3(n2591), .A4(n2590), .ZN(n2604)
         );
  OAI22_X1 U2656 ( .A1(n345), .A2(n3777), .B1(n665), .B2(n3756), .ZN(n2597) );
  OAI22_X1 U2657 ( .A1(n601), .A2(n3759), .B1(n313), .B2(n3764), .ZN(n2596) );
  OAI22_X1 U2658 ( .A1(n697), .A2(n3765), .B1(n537), .B2(n3779), .ZN(n2595) );
  OAI22_X1 U2659 ( .A1(n569), .A2(n3782), .B1(n121), .B2(n3774), .ZN(n2594) );
  NOR4_X1 U2660 ( .A1(n2597), .A2(n2596), .A3(n2595), .A4(n2594), .ZN(n2603)
         );
  OAI22_X1 U2661 ( .A1(n921), .A2(n3783), .B1(n633), .B2(n3755), .ZN(n2601) );
  OAI22_X1 U2662 ( .A1(n249), .A2(n3781), .B1(n793), .B2(n3772), .ZN(n2600) );
  OAI22_X1 U2663 ( .A1(n377), .A2(n3776), .B1(n857), .B2(n3767), .ZN(n2599) );
  OAI22_X1 U2664 ( .A1(n729), .A2(n3762), .B1(n505), .B2(n3757), .ZN(n2598) );
  NOR4_X1 U2665 ( .A1(n2601), .A2(n2600), .A3(n2599), .A4(n2598), .ZN(n2602)
         );
  NAND4_X1 U2666 ( .A1(n2605), .A2(n2604), .A3(n2603), .A4(n2602), .ZN(n2606)
         );
  AOI22_X1 U2667 ( .A1(lo_out[24]), .A2(n3786), .B1(n3785), .B2(n2606), .ZN(
        n2607) );
  OAI21_X1 U2668 ( .B1(n1642), .B2(n3787), .A(n2607), .ZN(rp2[24]) );
  NOR2_X1 U2669 ( .A1(n378), .A2(n3776), .ZN(n2611) );
  OAI22_X1 U2670 ( .A1(n602), .A2(n3759), .B1(n762), .B2(n3768), .ZN(n2610) );
  OAI22_X1 U2671 ( .A1(n218), .A2(n3758), .B1(n730), .B2(n3762), .ZN(n2609) );
  OAI22_X1 U2672 ( .A1(n698), .A2(n3765), .B1(n154), .B2(n1682), .ZN(n2608) );
  NOR4_X1 U2673 ( .A1(n2611), .A2(n2610), .A3(n2609), .A4(n2608), .ZN(n3619)
         );
  OAI22_X1 U2674 ( .A1(n474), .A2(n3766), .B1(n58), .B2(n3773), .ZN(n2615) );
  OAI22_X1 U2675 ( .A1(n410), .A2(n3780), .B1(n826), .B2(n3754), .ZN(n2614) );
  OAI22_X1 U2676 ( .A1(n666), .A2(n3756), .B1(n922), .B2(n3783), .ZN(n2613) );
  OAI22_X1 U2677 ( .A1(n314), .A2(n3764), .B1(n506), .B2(n3757), .ZN(n2612) );
  NOR4_X1 U2678 ( .A1(n2615), .A2(n2614), .A3(n2613), .A4(n2612), .ZN(n3618)
         );
  OAI22_X1 U2679 ( .A1(n954), .A2(n3784), .B1(n122), .B2(n3774), .ZN(n2619) );
  OAI22_X1 U2680 ( .A1(n346), .A2(n3777), .B1(n986), .B2(n3771), .ZN(n2618) );
  OAI22_X1 U2681 ( .A1(n634), .A2(n1681), .B1(n538), .B2(n3779), .ZN(n2617) );
  OAI22_X1 U2682 ( .A1(n90), .A2(n3763), .B1(n186), .B2(n3761), .ZN(n2616) );
  NOR4_X1 U2683 ( .A1(n2619), .A2(n2618), .A3(n2617), .A4(n2616), .ZN(n3617)
         );
  OAI22_X1 U2684 ( .A1(n858), .A2(n3767), .B1(n250), .B2(n3781), .ZN(n3615) );
  OAI22_X1 U2685 ( .A1(n26), .A2(n3770), .B1(n282), .B2(n3775), .ZN(n2622) );
  OAI22_X1 U2686 ( .A1(n570), .A2(n3782), .B1(n890), .B2(n3778), .ZN(n2621) );
  OAI22_X1 U2687 ( .A1(n794), .A2(n3772), .B1(n442), .B2(n3760), .ZN(n2620) );
  NOR4_X1 U2688 ( .A1(n3615), .A2(n2622), .A3(n2621), .A4(n2620), .ZN(n3616)
         );
  NAND4_X1 U2689 ( .A1(n3619), .A2(n3618), .A3(n3617), .A4(n3616), .ZN(n3620)
         );
  AOI22_X1 U2690 ( .A1(lo_out[25]), .A2(n3786), .B1(n1684), .B2(n3620), .ZN(
        n3621) );
  OAI21_X1 U2691 ( .B1(n1652), .B2(n3787), .A(n3621), .ZN(rp2[25]) );
  NOR2_X1 U2692 ( .A1(n795), .A2(n3772), .ZN(n3625) );
  OAI22_X1 U2693 ( .A1(n667), .A2(n3756), .B1(n731), .B2(n3762), .ZN(n3624) );
  OAI22_X1 U2694 ( .A1(n859), .A2(n3767), .B1(n827), .B2(n3754), .ZN(n3623) );
  OAI22_X1 U2695 ( .A1(n123), .A2(n3774), .B1(n59), .B2(n3773), .ZN(n3622) );
  NOR4_X1 U2696 ( .A1(n3625), .A2(n3624), .A3(n3623), .A4(n3622), .ZN(n3641)
         );
  OAI22_X1 U2697 ( .A1(n155), .A2(n1682), .B1(n635), .B2(n3755), .ZN(n3629) );
  OAI22_X1 U2698 ( .A1(n347), .A2(n3777), .B1(n379), .B2(n3776), .ZN(n3628) );
  OAI22_X1 U2699 ( .A1(n187), .A2(n3761), .B1(n891), .B2(n3778), .ZN(n3627) );
  OAI22_X1 U2700 ( .A1(n91), .A2(n3763), .B1(n443), .B2(n3760), .ZN(n3626) );
  NOR4_X1 U2701 ( .A1(n3629), .A2(n3628), .A3(n3627), .A4(n3626), .ZN(n3640)
         );
  OAI22_X1 U2702 ( .A1(n219), .A2(n3758), .B1(n539), .B2(n3779), .ZN(n3633) );
  OAI22_X1 U2703 ( .A1(n603), .A2(n3759), .B1(n283), .B2(n3775), .ZN(n3632) );
  OAI22_X1 U2704 ( .A1(n763), .A2(n3768), .B1(n955), .B2(n3784), .ZN(n3631) );
  OAI22_X1 U2705 ( .A1(n507), .A2(n3757), .B1(n923), .B2(n3783), .ZN(n3630) );
  NOR4_X1 U2706 ( .A1(n3633), .A2(n3632), .A3(n3631), .A4(n3630), .ZN(n3639)
         );
  OAI22_X1 U2707 ( .A1(n987), .A2(n3771), .B1(n315), .B2(n3764), .ZN(n3637) );
  OAI22_X1 U2708 ( .A1(n571), .A2(n3782), .B1(n699), .B2(n3765), .ZN(n3636) );
  OAI22_X1 U2709 ( .A1(n411), .A2(n3780), .B1(n475), .B2(n3766), .ZN(n3635) );
  OAI22_X1 U2710 ( .A1(n27), .A2(n3770), .B1(n251), .B2(n3781), .ZN(n3634) );
  NOR4_X1 U2711 ( .A1(n3637), .A2(n3636), .A3(n3635), .A4(n3634), .ZN(n3638)
         );
  NAND4_X1 U2712 ( .A1(n3641), .A2(n3640), .A3(n3639), .A4(n3638), .ZN(n3642)
         );
  AOI22_X1 U2713 ( .A1(lo_out[26]), .A2(n1685), .B1(n1684), .B2(n3642), .ZN(
        n3643) );
  OAI21_X1 U2714 ( .B1(n1643), .B2(n3787), .A(n3643), .ZN(rp2[26]) );
  NOR2_X1 U2715 ( .A1(n252), .A2(n3781), .ZN(n3647) );
  OAI22_X1 U2716 ( .A1(n92), .A2(n3763), .B1(n732), .B2(n3762), .ZN(n3646) );
  OAI22_X1 U2717 ( .A1(n828), .A2(n3754), .B1(n540), .B2(n3779), .ZN(n3645) );
  OAI22_X1 U2718 ( .A1(n700), .A2(n3765), .B1(n796), .B2(n3772), .ZN(n3644) );
  NOR4_X1 U2719 ( .A1(n3647), .A2(n3646), .A3(n3645), .A4(n3644), .ZN(n3663)
         );
  OAI22_X1 U2720 ( .A1(n188), .A2(n3761), .B1(n156), .B2(n1682), .ZN(n3651) );
  OAI22_X1 U2721 ( .A1(n412), .A2(n3780), .B1(n476), .B2(n3766), .ZN(n3650) );
  OAI22_X1 U2722 ( .A1(n28), .A2(n3770), .B1(n284), .B2(n3775), .ZN(n3649) );
  OAI22_X1 U2723 ( .A1(n572), .A2(n3782), .B1(n444), .B2(n3760), .ZN(n3648) );
  NOR4_X1 U2724 ( .A1(n3651), .A2(n3650), .A3(n3649), .A4(n3648), .ZN(n3662)
         );
  OAI22_X1 U2725 ( .A1(n380), .A2(n3776), .B1(n508), .B2(n3757), .ZN(n3655) );
  OAI22_X1 U2726 ( .A1(n892), .A2(n3778), .B1(n860), .B2(n3767), .ZN(n3654) );
  OAI22_X1 U2727 ( .A1(n220), .A2(n3758), .B1(n924), .B2(n3783), .ZN(n3653) );
  OAI22_X1 U2728 ( .A1(n636), .A2(n1681), .B1(n348), .B2(n3777), .ZN(n3652) );
  NOR4_X1 U2729 ( .A1(n3655), .A2(n3654), .A3(n3653), .A4(n3652), .ZN(n3661)
         );
  OAI22_X1 U2730 ( .A1(n956), .A2(n3784), .B1(n124), .B2(n3774), .ZN(n3659) );
  OAI22_X1 U2731 ( .A1(n316), .A2(n3764), .B1(n988), .B2(n3771), .ZN(n3658) );
  OAI22_X1 U2732 ( .A1(n668), .A2(n3756), .B1(n60), .B2(n3773), .ZN(n3657) );
  OAI22_X1 U2733 ( .A1(n764), .A2(n3768), .B1(n604), .B2(n3759), .ZN(n3656) );
  NOR4_X1 U2734 ( .A1(n3659), .A2(n3658), .A3(n3657), .A4(n3656), .ZN(n3660)
         );
  NAND4_X1 U2735 ( .A1(n3663), .A2(n3662), .A3(n3661), .A4(n3660), .ZN(n3664)
         );
  AOI22_X1 U2736 ( .A1(lo_out[27]), .A2(n1685), .B1(n3785), .B2(n3664), .ZN(
        n3665) );
  OAI21_X1 U2737 ( .B1(n1644), .B2(n3787), .A(n3665), .ZN(rp2[27]) );
  NOR2_X1 U2738 ( .A1(n509), .A2(n3757), .ZN(n3669) );
  OAI22_X1 U2739 ( .A1(n61), .A2(n3773), .B1(n765), .B2(n3768), .ZN(n3668) );
  OAI22_X1 U2740 ( .A1(n861), .A2(n3767), .B1(n701), .B2(n3765), .ZN(n3667) );
  OAI22_X1 U2741 ( .A1(n381), .A2(n3776), .B1(n797), .B2(n3772), .ZN(n3666) );
  NOR4_X1 U2742 ( .A1(n3669), .A2(n3668), .A3(n3667), .A4(n3666), .ZN(n3685)
         );
  OAI22_X1 U2743 ( .A1(n477), .A2(n3766), .B1(n285), .B2(n3775), .ZN(n3673) );
  OAI22_X1 U2744 ( .A1(n733), .A2(n3762), .B1(n221), .B2(n3758), .ZN(n3672) );
  OAI22_X1 U2745 ( .A1(n253), .A2(n3781), .B1(n605), .B2(n3759), .ZN(n3671) );
  OAI22_X1 U2746 ( .A1(n957), .A2(n3784), .B1(n541), .B2(n3779), .ZN(n3670) );
  NOR4_X1 U2747 ( .A1(n3673), .A2(n3672), .A3(n3671), .A4(n3670), .ZN(n3684)
         );
  OAI22_X1 U2748 ( .A1(n989), .A2(n3771), .B1(n93), .B2(n3763), .ZN(n3677) );
  OAI22_X1 U2749 ( .A1(n29), .A2(n3770), .B1(n669), .B2(n3756), .ZN(n3676) );
  OAI22_X1 U2750 ( .A1(n125), .A2(n3774), .B1(n157), .B2(n3769), .ZN(n3675) );
  OAI22_X1 U2751 ( .A1(n349), .A2(n3777), .B1(n317), .B2(n3764), .ZN(n3674) );
  NOR4_X1 U2752 ( .A1(n3677), .A2(n3676), .A3(n3675), .A4(n3674), .ZN(n3683)
         );
  OAI22_X1 U2753 ( .A1(n189), .A2(n3761), .B1(n925), .B2(n3783), .ZN(n3681) );
  OAI22_X1 U2754 ( .A1(n445), .A2(n3760), .B1(n829), .B2(n3754), .ZN(n3680) );
  OAI22_X1 U2755 ( .A1(n893), .A2(n3778), .B1(n573), .B2(n3782), .ZN(n3679) );
  OAI22_X1 U2756 ( .A1(n413), .A2(n3780), .B1(n637), .B2(n3755), .ZN(n3678) );
  NOR4_X1 U2757 ( .A1(n3681), .A2(n3680), .A3(n3679), .A4(n3678), .ZN(n3682)
         );
  NAND4_X1 U2758 ( .A1(n3685), .A2(n3684), .A3(n3683), .A4(n3682), .ZN(n3686)
         );
  AOI22_X1 U2759 ( .A1(lo_out[28]), .A2(n1685), .B1(n3785), .B2(n3686), .ZN(
        n3687) );
  OAI21_X1 U2760 ( .B1(n1645), .B2(n3787), .A(n3687), .ZN(rp2[28]) );
  NOR2_X1 U2761 ( .A1(n222), .A2(n3758), .ZN(n3691) );
  OAI22_X1 U2762 ( .A1(n670), .A2(n3756), .B1(n62), .B2(n3773), .ZN(n3690) );
  OAI22_X1 U2763 ( .A1(n702), .A2(n3765), .B1(n638), .B2(n3755), .ZN(n3689) );
  OAI22_X1 U2764 ( .A1(n766), .A2(n3768), .B1(n830), .B2(n3754), .ZN(n3688) );
  NOR4_X1 U2765 ( .A1(n3691), .A2(n3690), .A3(n3689), .A4(n3688), .ZN(n3707)
         );
  OAI22_X1 U2766 ( .A1(n862), .A2(n3767), .B1(n734), .B2(n3762), .ZN(n3695) );
  OAI22_X1 U2767 ( .A1(n990), .A2(n3771), .B1(n510), .B2(n3757), .ZN(n3694) );
  OAI22_X1 U2768 ( .A1(n894), .A2(n3778), .B1(n318), .B2(n3764), .ZN(n3693) );
  OAI22_X1 U2769 ( .A1(n446), .A2(n3760), .B1(n94), .B2(n3763), .ZN(n3692) );
  NOR4_X1 U2770 ( .A1(n3695), .A2(n3694), .A3(n3693), .A4(n3692), .ZN(n3706)
         );
  OAI22_X1 U2771 ( .A1(n158), .A2(n1682), .B1(n382), .B2(n3776), .ZN(n3699) );
  OAI22_X1 U2772 ( .A1(n606), .A2(n3759), .B1(n286), .B2(n3775), .ZN(n3698) );
  OAI22_X1 U2773 ( .A1(n190), .A2(n3761), .B1(n926), .B2(n3783), .ZN(n3697) );
  OAI22_X1 U2774 ( .A1(n574), .A2(n3782), .B1(n958), .B2(n3784), .ZN(n3696) );
  NOR4_X1 U2775 ( .A1(n3699), .A2(n3698), .A3(n3697), .A4(n3696), .ZN(n3705)
         );
  OAI22_X1 U2776 ( .A1(n30), .A2(n3770), .B1(n126), .B2(n3774), .ZN(n3703) );
  OAI22_X1 U2777 ( .A1(n542), .A2(n3779), .B1(n478), .B2(n3766), .ZN(n3702) );
  OAI22_X1 U2778 ( .A1(n254), .A2(n3781), .B1(n350), .B2(n3777), .ZN(n3701) );
  OAI22_X1 U2779 ( .A1(n414), .A2(n3780), .B1(n798), .B2(n3772), .ZN(n3700) );
  NOR4_X1 U2780 ( .A1(n3703), .A2(n3702), .A3(n3701), .A4(n3700), .ZN(n3704)
         );
  NAND4_X1 U2781 ( .A1(n3707), .A2(n3706), .A3(n3705), .A4(n3704), .ZN(n3708)
         );
  AOI22_X1 U2782 ( .A1(lo_out[29]), .A2(n1685), .B1(n1684), .B2(n3708), .ZN(
        n3709) );
  OAI21_X1 U2783 ( .B1(n1646), .B2(n3787), .A(n3709), .ZN(rp2[29]) );
  NOR2_X1 U2784 ( .A1(n351), .A2(n3777), .ZN(n3713) );
  OAI22_X1 U2785 ( .A1(n319), .A2(n3764), .B1(n767), .B2(n3768), .ZN(n3712) );
  OAI22_X1 U2786 ( .A1(n95), .A2(n3763), .B1(n735), .B2(n3762), .ZN(n3711) );
  OAI22_X1 U2787 ( .A1(n895), .A2(n3778), .B1(n959), .B2(n3784), .ZN(n3710) );
  NOR4_X1 U2788 ( .A1(n3713), .A2(n3712), .A3(n3711), .A4(n3710), .ZN(n3729)
         );
  OAI22_X1 U2789 ( .A1(n159), .A2(n1682), .B1(n479), .B2(n3766), .ZN(n3717) );
  OAI22_X1 U2790 ( .A1(n543), .A2(n3779), .B1(n831), .B2(n3754), .ZN(n3716) );
  OAI22_X1 U2791 ( .A1(n703), .A2(n3765), .B1(n927), .B2(n3783), .ZN(n3715) );
  OAI22_X1 U2792 ( .A1(n287), .A2(n3775), .B1(n63), .B2(n3773), .ZN(n3714) );
  NOR4_X1 U2793 ( .A1(n3717), .A2(n3716), .A3(n3715), .A4(n3714), .ZN(n3728)
         );
  OAI22_X1 U2794 ( .A1(n607), .A2(n3759), .B1(n575), .B2(n3782), .ZN(n3721) );
  OAI22_X1 U2795 ( .A1(n863), .A2(n3767), .B1(n223), .B2(n3758), .ZN(n3720) );
  OAI22_X1 U2796 ( .A1(n255), .A2(n3781), .B1(n799), .B2(n3772), .ZN(n3719) );
  OAI22_X1 U2797 ( .A1(n383), .A2(n3776), .B1(n639), .B2(n3755), .ZN(n3718) );
  NOR4_X1 U2798 ( .A1(n3721), .A2(n3720), .A3(n3719), .A4(n3718), .ZN(n3727)
         );
  OAI22_X1 U2799 ( .A1(n191), .A2(n3761), .B1(n127), .B2(n3774), .ZN(n3725) );
  OAI22_X1 U2800 ( .A1(n415), .A2(n3780), .B1(n511), .B2(n3757), .ZN(n3724) );
  OAI22_X1 U2801 ( .A1(n31), .A2(n3770), .B1(n671), .B2(n3756), .ZN(n3723) );
  OAI22_X1 U2802 ( .A1(n991), .A2(n3771), .B1(n447), .B2(n3760), .ZN(n3722) );
  NOR4_X1 U2803 ( .A1(n3725), .A2(n3724), .A3(n3723), .A4(n3722), .ZN(n3726)
         );
  NAND4_X1 U2804 ( .A1(n3729), .A2(n3728), .A3(n3727), .A4(n3726), .ZN(n3730)
         );
  AOI22_X1 U2805 ( .A1(lo_out[30]), .A2(n1685), .B1(n3785), .B2(n3730), .ZN(
        n3731) );
  OAI21_X1 U2806 ( .B1(n1654), .B2(n3787), .A(n3731), .ZN(rp2[30]) );
  NOR2_X1 U2807 ( .A1(n960), .A2(n3784), .ZN(n3735) );
  OAI22_X1 U2808 ( .A1(n64), .A2(n3773), .B1(n288), .B2(n3775), .ZN(n3734) );
  OAI22_X1 U2809 ( .A1(n640), .A2(n3755), .B1(n320), .B2(n3764), .ZN(n3733) );
  OAI22_X1 U2810 ( .A1(n576), .A2(n3782), .B1(n96), .B2(n3763), .ZN(n3732) );
  NOR4_X1 U2811 ( .A1(n3735), .A2(n3734), .A3(n3733), .A4(n3732), .ZN(n3751)
         );
  OAI22_X1 U2812 ( .A1(n608), .A2(n3759), .B1(n192), .B2(n3761), .ZN(n3739) );
  OAI22_X1 U2813 ( .A1(n32), .A2(n3770), .B1(n352), .B2(n3777), .ZN(n3738) );
  OAI22_X1 U2814 ( .A1(n992), .A2(n3771), .B1(n128), .B2(n3774), .ZN(n3737) );
  OAI22_X1 U2815 ( .A1(n800), .A2(n3772), .B1(n480), .B2(n3766), .ZN(n3736) );
  NOR4_X1 U2816 ( .A1(n3739), .A2(n3738), .A3(n3737), .A4(n3736), .ZN(n3750)
         );
  OAI22_X1 U2817 ( .A1(n928), .A2(n3783), .B1(n160), .B2(n1682), .ZN(n3743) );
  OAI22_X1 U2818 ( .A1(n416), .A2(n3780), .B1(n768), .B2(n3768), .ZN(n3742) );
  OAI22_X1 U2819 ( .A1(n224), .A2(n3758), .B1(n864), .B2(n3767), .ZN(n3741) );
  OAI22_X1 U2820 ( .A1(n672), .A2(n3756), .B1(n736), .B2(n3762), .ZN(n3740) );
  NOR4_X1 U2821 ( .A1(n3743), .A2(n3742), .A3(n3741), .A4(n3740), .ZN(n3749)
         );
  OAI22_X1 U2822 ( .A1(n512), .A2(n3757), .B1(n704), .B2(n3765), .ZN(n3747) );
  OAI22_X1 U2823 ( .A1(n896), .A2(n3778), .B1(n544), .B2(n3779), .ZN(n3746) );
  OAI22_X1 U2824 ( .A1(n448), .A2(n3760), .B1(n256), .B2(n3781), .ZN(n3745) );
  OAI22_X1 U2825 ( .A1(n832), .A2(n3754), .B1(n384), .B2(n3776), .ZN(n3744) );
  NOR4_X1 U2826 ( .A1(n3747), .A2(n3746), .A3(n3745), .A4(n3744), .ZN(n3748)
         );
  NAND4_X1 U2827 ( .A1(n3751), .A2(n3750), .A3(n3749), .A4(n3748), .ZN(n3752)
         );
  AOI22_X1 U2828 ( .A1(lo_out[31]), .A2(n3786), .B1(n1684), .B2(n3752), .ZN(
        n3753) );
  OAI21_X1 U2829 ( .B1(n1647), .B2(n3787), .A(n3753), .ZN(rp2[31]) );
endmodule


module shifter_t2 ( data_in, shift, shift_type, data_out );
  input [31:0] data_in;
  input [4:0] shift;
  input [3:0] shift_type;
  output [31:0] data_out;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834;

  OAI33_X1 U2 ( .A1(1'b0), .A2(n138), .A3(n52), .B1(n62), .B2(n673), .B3(n129), 
        .ZN(n123) );
  INV_X2 U3 ( .A(n795), .ZN(n792) );
  AOI211_X1 U4 ( .C1(n784), .C2(n613), .A(n612), .B(n611), .ZN(n1) );
  NAND4_X1 U5 ( .A1(n642), .A2(n643), .A3(n1), .A4(n644), .ZN(data_out[31]) );
  OAI211_X1 U6 ( .C1(n531), .C2(n827), .A(n530), .B(n529), .ZN(data_out[29])
         );
  AOI22_X1 U7 ( .A1(n568), .A2(n132), .B1(n502), .B2(n138), .ZN(n2) );
  AOI22_X1 U8 ( .A1(n295), .A2(n175), .B1(n551), .B2(n183), .ZN(n3) );
  OAI22_X1 U9 ( .A1(n708), .A2(n668), .B1(n683), .B2(n834), .ZN(n4) );
  OAI22_X1 U10 ( .A1(n134), .A2(n652), .B1(n135), .B2(n651), .ZN(n5) );
  OAI22_X1 U11 ( .A1(n628), .A2(n137), .B1(n142), .B2(n136), .ZN(n6) );
  OR4_X1 U12 ( .A1(n800), .A2(n4), .A3(n5), .A4(n6), .ZN(n7) );
  AOI221_X1 U13 ( .B1(n143), .B2(n258), .C1(n164), .C2(n258), .A(n7), .ZN(n8)
         );
  OAI21_X1 U14 ( .B1(n170), .B2(n153), .A(n553), .ZN(n9) );
  NAND4_X1 U15 ( .A1(n2), .A2(n3), .A3(n8), .A4(n9), .ZN(data_out[12]) );
  OAI22_X1 U16 ( .A1(n585), .A2(n816), .B1(n474), .B2(n834), .ZN(n10) );
  OAI211_X1 U17 ( .C1(n629), .C2(n668), .A(n644), .B(n504), .ZN(n11) );
  AOI211_X1 U18 ( .C1(n443), .C2(n619), .A(n10), .B(n11), .ZN(n12) );
  OAI22_X1 U19 ( .A1(n506), .A2(n709), .B1(n444), .B2(n660), .ZN(n13) );
  OAI22_X1 U20 ( .A1(n628), .A2(n467), .B1(n579), .B2(n678), .ZN(n14) );
  NOR3_X1 U21 ( .A1(n465), .A2(n13), .A3(n14), .ZN(n15) );
  OAI211_X1 U22 ( .C1(n472), .C2(n614), .A(n12), .B(n15), .ZN(data_out[27]) );
  AOI22_X1 U23 ( .A1(n339), .A2(n502), .B1(n618), .B2(n634), .ZN(n16) );
  OAI22_X1 U24 ( .A1(n797), .A2(n354), .B1(n827), .B2(n326), .ZN(n17) );
  OAI22_X1 U25 ( .A1(n378), .A2(n719), .B1(n327), .B2(n660), .ZN(n18) );
  OAI22_X1 U26 ( .A1(n379), .A2(n709), .B1(n328), .B2(n651), .ZN(n19) );
  AOI211_X1 U27 ( .C1(n564), .C2(n632), .A(n336), .B(n335), .ZN(n20) );
  OAI21_X1 U28 ( .B1(n816), .B2(n342), .A(n20), .ZN(n21) );
  NOR4_X1 U29 ( .A1(n17), .A2(n18), .A3(n19), .A4(n21), .ZN(n22) );
  OAI211_X1 U30 ( .C1(n637), .C2(n337), .A(n16), .B(n22), .ZN(data_out[22]) );
  OAI22_X1 U31 ( .A1(n481), .A2(n364), .B1(n193), .B2(n605), .ZN(n23) );
  AOI221_X1 U32 ( .B1(n194), .B2(n551), .C1(n254), .C2(n551), .A(n23), .ZN(n24) );
  OAI21_X1 U33 ( .B1(n219), .B2(n234), .A(n258), .ZN(n25) );
  OAI21_X1 U34 ( .B1(n200), .B2(n250), .A(n295), .ZN(n26) );
  OAI21_X1 U35 ( .B1(n240), .B2(n213), .A(n553), .ZN(n27) );
  NAND4_X1 U36 ( .A1(n24), .A2(n25), .A3(n26), .A4(n27), .ZN(data_out[16]) );
  INV_X1 U37 ( .A(n652), .ZN(n28) );
  AOI22_X1 U38 ( .A1(n295), .A2(n164), .B1(n116), .B2(n28), .ZN(n29) );
  OAI21_X1 U39 ( .B1(n112), .B2(n136), .A(n824), .ZN(n30) );
  OAI22_X1 U40 ( .A1(n683), .A2(n668), .B1(n142), .B2(n625), .ZN(n31) );
  AOI211_X1 U41 ( .C1(n114), .C2(n778), .A(n30), .B(n31), .ZN(n32) );
  INV_X1 U42 ( .A(n170), .ZN(n33) );
  OAI22_X1 U43 ( .A1(n715), .A2(n33), .B1(n123), .B2(n812), .ZN(n34) );
  AOI22_X1 U44 ( .A1(n132), .A2(n502), .B1(n658), .B2(n802), .ZN(n35) );
  OAI21_X1 U45 ( .B1(n628), .B2(n135), .A(n35), .ZN(n36) );
  AOI211_X1 U46 ( .C1(n553), .C2(n143), .A(n34), .B(n36), .ZN(n37) );
  AOI22_X1 U47 ( .A1(n258), .A2(n153), .B1(n117), .B2(n118), .ZN(n38) );
  NAND4_X1 U48 ( .A1(n29), .A2(n32), .A3(n37), .A4(n38), .ZN(data_out[11]) );
  AOI22_X1 U49 ( .A1(n778), .A2(n809), .B1(n114), .B2(n810), .ZN(n39) );
  AOI22_X1 U50 ( .A1(n551), .A2(n143), .B1(n802), .B2(n822), .ZN(n40) );
  AOI22_X1 U51 ( .A1(n808), .A2(n563), .B1(n658), .B2(n823), .ZN(n41) );
  OAI22_X1 U52 ( .A1(n818), .A2(n123), .B1(n812), .B2(n819), .ZN(n42) );
  AOI22_X1 U53 ( .A1(n821), .A2(n815), .B1(n116), .B2(n118), .ZN(n43) );
  OAI211_X1 U54 ( .C1(n112), .C2(n625), .A(n824), .B(n43), .ZN(n44) );
  AOI211_X1 U55 ( .C1(n295), .C2(n153), .A(n42), .B(n44), .ZN(n45) );
  NAND4_X1 U56 ( .A1(n39), .A2(n40), .A3(n41), .A4(n45), .ZN(data_out[10]) );
  AOI22_X1 U57 ( .A1(n802), .A2(n820), .B1(n823), .B2(n544), .ZN(n46) );
  AOI22_X1 U58 ( .A1(n551), .A2(n552), .B1(n778), .B2(n266), .ZN(n47) );
  AOI22_X1 U59 ( .A1(n822), .A2(n765), .B1(n775), .B2(n740), .ZN(n48) );
  OAI22_X1 U60 ( .A1(n718), .A2(n670), .B1(n812), .B2(n271), .ZN(n49) );
  OAI22_X1 U61 ( .A1(n547), .A2(n549), .B1(n548), .B2(n545), .ZN(n50) );
  AOI211_X1 U62 ( .C1(n821), .C2(n272), .A(n49), .B(n50), .ZN(n51) );
  NAND4_X1 U63 ( .A1(n46), .A2(n47), .A3(n48), .A4(n51), .ZN(data_out[1]) );
  INV_X1 U64 ( .A(n62), .ZN(n52) );
  OAI21_X1 U66 ( .B1(n219), .B2(n164), .A(n551), .ZN(n54) );
  OAI21_X1 U67 ( .B1(n768), .B2(n668), .A(n54), .ZN(n55) );
  AOI211_X1 U68 ( .C1(n741), .C2(n802), .A(n800), .B(n55), .ZN(n56) );
  OAI21_X1 U69 ( .B1(n175), .B2(n200), .A(n553), .ZN(n57) );
  OAI21_X1 U70 ( .B1(n213), .B2(n170), .A(n295), .ZN(n58) );
  OAI21_X1 U71 ( .B1(n194), .B2(n183), .A(n258), .ZN(n59) );
  NAND4_X1 U72 ( .A1(n56), .A2(n57), .A3(n58), .A4(n59), .ZN(data_out[14]) );
  INV_X1 U73 ( .A(n62), .ZN(n60) );
  NAND2_X1 U74 ( .A1(n696), .A2(n60), .ZN(n61) );
  OAI22_X1 U75 ( .A1(n121), .A2(n61), .B1(n132), .B2(n60), .ZN(n819) );
  INV_X2 U76 ( .A(n604), .ZN(n607) );
  INV_X2 U77 ( .A(shift[2]), .ZN(n70) );
  INV_X2 U78 ( .A(n760), .ZN(n789) );
  INV_X4 U79 ( .A(n70), .ZN(n63) );
  INV_X2 U80 ( .A(n758), .ZN(n787) );
  INV_X1 U81 ( .A(n757), .ZN(n786) );
  AND3_X1 U82 ( .A1(n65), .A2(n66), .A3(data_in[31]), .ZN(n64) );
  INV_X1 U83 ( .A(n834), .ZN(n802) );
  INV_X1 U84 ( .A(n669), .ZN(n553) );
  INV_X1 U85 ( .A(n668), .ZN(n823) );
  INV_X1 U86 ( .A(n69), .ZN(n67) );
  INV_X2 U87 ( .A(n71), .ZN(n62) );
  INV_X1 U88 ( .A(shift[0]), .ZN(n400) );
  OAI22_X4 U89 ( .A1(n74), .A2(shift_type[0]), .B1(n101), .B2(shift_type[0]), 
        .ZN(n533) );
  OR4_X1 U90 ( .A1(n695), .A2(n694), .A3(n693), .A4(n692), .ZN(data_out[4]) );
  NOR2_X1 U91 ( .A1(n67), .A2(n264), .ZN(n681) );
  INV_X1 U92 ( .A(n340), .ZN(n333) );
  INV_X1 U93 ( .A(n111), .ZN(n297) );
  INV_X1 U94 ( .A(n535), .ZN(n536) );
  INV_X1 U95 ( .A(n69), .ZN(n68) );
  NAND2_X1 U96 ( .A1(n72), .A2(n70), .ZN(n758) );
  NAND2_X1 U97 ( .A1(n70), .A2(n62), .ZN(n795) );
  NAND2_X1 U98 ( .A1(n72), .A2(n63), .ZN(n760) );
  NAND2_X1 U99 ( .A1(n62), .A2(n63), .ZN(n757) );
  INV_X1 U100 ( .A(shift[1]), .ZN(n72) );
  INV_X1 U101 ( .A(n64), .ZN(n605) );
  INV_X1 U102 ( .A(n534), .ZN(n537) );
  INV_X1 U103 ( .A(n671), .ZN(n258) );
  INV_X1 U104 ( .A(shift[1]), .ZN(n71) );
  BUF_X2 U105 ( .A(n70), .Z(n69) );
  INV_X1 U106 ( .A(n348), .ZN(n366) );
  NOR2_X2 U107 ( .A1(n71), .A2(n400), .ZN(n295) );
  NOR2_X2 U108 ( .A1(n62), .A2(shift[0]), .ZN(n551) );
  NOR3_X2 U109 ( .A1(n66), .A2(shift[3]), .A3(shift[4]), .ZN(n265) );
  INV_X1 U110 ( .A(n481), .ZN(n634) );
  NAND2_X1 U111 ( .A1(n80), .A2(n100), .ZN(n535) );
  INV_X1 U112 ( .A(n523), .ZN(n632) );
  INV_X1 U113 ( .A(n101), .ZN(n65) );
  NAND2_X1 U114 ( .A1(shift[3]), .A2(n80), .ZN(n534) );
  INV_X1 U115 ( .A(shift_type[2]), .ZN(n75) );
  INV_X1 U116 ( .A(shift_type[0]), .ZN(n66) );
  NOR2_X1 U117 ( .A1(shift_type[0]), .A2(shift[4]), .ZN(n80) );
  INV_X1 U118 ( .A(shift[3]), .ZN(n100) );
  NOR2_X1 U119 ( .A1(n400), .A2(n535), .ZN(n782) );
  INV_X1 U120 ( .A(n782), .ZN(n818) );
  INV_X1 U121 ( .A(shift_type[1]), .ZN(n73) );
  OR2_X1 U122 ( .A1(n73), .A2(shift_type[2]), .ZN(n74) );
  NAND2_X1 U123 ( .A1(shift_type[2]), .A2(n73), .ZN(n101) );
  INV_X1 U124 ( .A(n533), .ZN(n264) );
  NAND3_X1 U125 ( .A1(shift_type[0]), .A2(shift_type[1]), .A3(n75), .ZN(n604)
         );
  NAND2_X1 U126 ( .A1(n607), .A2(data_in[0]), .ZN(n283) );
  INV_X1 U127 ( .A(n283), .ZN(n320) );
  NOR2_X1 U128 ( .A1(n69), .A2(n264), .ZN(n88) );
  AOI22_X1 U129 ( .A1(n68), .A2(n320), .B1(data_in[7]), .B2(n88), .ZN(n76) );
  INV_X1 U130 ( .A(n76), .ZN(n672) );
  AOI21_X1 U131 ( .B1(data_in[3]), .B2(n681), .A(n672), .ZN(n661) );
  INV_X1 U132 ( .A(data_in[5]), .ZN(n305) );
  AOI22_X1 U133 ( .A1(n62), .A2(n661), .B1(n789), .B2(n305), .ZN(n77) );
  OAI211_X1 U134 ( .C1(data_in[1]), .C2(n758), .A(n533), .B(n77), .ZN(n271) );
  INV_X1 U135 ( .A(shift[4]), .ZN(n192) );
  NOR2_X1 U136 ( .A1(n192), .A2(shift_type[0]), .ZN(n203) );
  NAND3_X1 U137 ( .A1(n100), .A2(shift[0]), .A3(n203), .ZN(n668) );
  NAND2_X1 U138 ( .A1(n533), .A2(data_in[21]), .ZN(n727) );
  INV_X1 U139 ( .A(data_in[23]), .ZN(n347) );
  INV_X1 U140 ( .A(n88), .ZN(n78) );
  NAND3_X1 U141 ( .A1(n533), .A2(data_in[19]), .A3(n69), .ZN(n128) );
  OAI21_X1 U142 ( .B1(n347), .B2(n78), .A(n128), .ZN(n116) );
  INV_X1 U143 ( .A(n116), .ZN(n543) );
  NAND2_X1 U144 ( .A1(n533), .A2(data_in[17]), .ZN(n729) );
  AOI222_X1 U145 ( .A1(n727), .A2(n789), .B1(n62), .B2(n543), .C1(n729), .C2(
        n787), .ZN(n820) );
  AOI22_X1 U146 ( .A1(data_in[15]), .A2(n88), .B1(data_in[11]), .B2(n681), 
        .ZN(n653) );
  OAI22_X1 U147 ( .A1(data_in[13]), .A2(n760), .B1(data_in[9]), .B2(n758), 
        .ZN(n79) );
  AOI211_X1 U148 ( .C1(n62), .C2(n653), .A(n264), .B(n79), .ZN(n272) );
  NOR2_X1 U149 ( .A1(n400), .A2(n534), .ZN(n776) );
  AOI22_X1 U150 ( .A1(n823), .A2(n820), .B1(n272), .B2(n776), .ZN(n97) );
  INV_X1 U151 ( .A(n203), .ZN(n193) );
  NOR2_X1 U152 ( .A1(shift[3]), .A2(n193), .ZN(n81) );
  NAND2_X1 U153 ( .A1(n81), .A2(n400), .ZN(n834) );
  NAND2_X1 U154 ( .A1(n533), .A2(data_in[16]), .ZN(n697) );
  INV_X1 U155 ( .A(n697), .ZN(n99) );
  INV_X1 U156 ( .A(data_in[22]), .ZN(n576) );
  NOR2_X1 U157 ( .A1(n264), .A2(n576), .ZN(n705) );
  OAI22_X1 U158 ( .A1(n99), .A2(n758), .B1(n705), .B2(n757), .ZN(n83) );
  NAND2_X1 U159 ( .A1(n533), .A2(data_in[20]), .ZN(n699) );
  INV_X1 U160 ( .A(n699), .ZN(n646) );
  NAND2_X1 U161 ( .A1(n533), .A2(data_in[18]), .ZN(n120) );
  INV_X1 U162 ( .A(n120), .ZN(n109) );
  OAI22_X1 U163 ( .A1(n646), .A2(n760), .B1(n109), .B2(n795), .ZN(n82) );
  NOR2_X1 U164 ( .A1(n83), .A2(n82), .ZN(n774) );
  AOI22_X1 U165 ( .A1(data_in[14]), .A2(n88), .B1(n681), .B2(data_in[10]), 
        .ZN(n548) );
  NAND2_X1 U166 ( .A1(n400), .A2(n62), .ZN(n671) );
  NAND2_X1 U167 ( .A1(n537), .A2(n258), .ZN(n684) );
  AOI22_X1 U168 ( .A1(n681), .A2(data_in[2]), .B1(data_in[6]), .B2(n88), .ZN(
        n549) );
  NOR2_X1 U169 ( .A1(n535), .A2(n671), .ZN(n493) );
  INV_X1 U170 ( .A(n493), .ZN(n719) );
  OAI22_X1 U171 ( .A1(n548), .A2(n684), .B1(n549), .B2(n719), .ZN(n95) );
  NAND2_X1 U172 ( .A1(n533), .A2(data_in[29]), .ZN(n331) );
  NAND2_X1 U173 ( .A1(n533), .A2(data_in[27]), .ZN(n124) );
  INV_X1 U174 ( .A(n124), .ZN(n195) );
  INV_X1 U175 ( .A(data_in[31]), .ZN(n606) );
  NOR2_X1 U176 ( .A1(n264), .A2(n606), .ZN(n365) );
  INV_X1 U177 ( .A(n365), .ZN(n188) );
  NAND2_X1 U178 ( .A1(n533), .A2(data_in[25]), .ZN(n104) );
  AOI22_X1 U179 ( .A1(n786), .A2(n188), .B1(n787), .B2(n104), .ZN(n84) );
  OAI21_X1 U180 ( .B1(n195), .B2(n795), .A(n84), .ZN(n85) );
  AOI21_X1 U181 ( .B1(n789), .B2(n331), .A(n85), .ZN(n775) );
  INV_X1 U182 ( .A(n775), .ZN(n833) );
  NAND2_X1 U183 ( .A1(shift[3]), .A2(n203), .ZN(n110) );
  NOR2_X1 U184 ( .A1(n400), .A2(n110), .ZN(n765) );
  INV_X1 U185 ( .A(n765), .ZN(n743) );
  INV_X1 U186 ( .A(data_in[8]), .ZN(n375) );
  NOR2_X1 U187 ( .A1(n535), .A2(shift[0]), .ZN(n784) );
  NAND2_X1 U188 ( .A1(data_in[0]), .A2(n784), .ZN(n86) );
  NAND2_X1 U189 ( .A1(n400), .A2(n537), .ZN(n637) );
  AOI221_X1 U190 ( .B1(n375), .B2(n86), .C1(n637), .C2(n86), .A(n758), .ZN(n89) );
  INV_X1 U191 ( .A(data_in[12]), .ZN(n268) );
  NAND2_X1 U192 ( .A1(n537), .A2(n551), .ZN(n652) );
  INV_X1 U193 ( .A(data_in[4]), .ZN(n267) );
  NAND2_X1 U194 ( .A1(n536), .A2(n551), .ZN(n660) );
  OAI22_X1 U195 ( .A1(n268), .A2(n652), .B1(n267), .B2(n660), .ZN(n87) );
  AOI22_X1 U196 ( .A1(n533), .A2(n89), .B1(n88), .B2(n87), .ZN(n93) );
  NAND2_X1 U197 ( .A1(n400), .A2(n265), .ZN(n798) );
  INV_X1 U198 ( .A(n798), .ZN(n810) );
  NOR2_X1 U199 ( .A1(n283), .A2(n63), .ZN(n796) );
  AOI21_X1 U200 ( .B1(n681), .B2(data_in[7]), .A(n796), .ZN(n674) );
  NOR2_X1 U201 ( .A1(n62), .A2(n674), .ZN(n266) );
  NOR2_X1 U202 ( .A1(shift[0]), .A2(n110), .ZN(n740) );
  INV_X1 U203 ( .A(data_in[28]), .ZN(n469) );
  NOR2_X1 U204 ( .A1(n264), .A2(n469), .ZN(n147) );
  INV_X1 U205 ( .A(n147), .ZN(n703) );
  NAND2_X1 U206 ( .A1(n533), .A2(data_in[26]), .ZN(n707) );
  INV_X1 U207 ( .A(n707), .ZN(n645) );
  NAND2_X1 U208 ( .A1(n533), .A2(data_in[30]), .ZN(n349) );
  NAND2_X1 U209 ( .A1(n533), .A2(data_in[24]), .ZN(n702) );
  AOI22_X1 U210 ( .A1(n786), .A2(n349), .B1(n787), .B2(n702), .ZN(n90) );
  OAI21_X1 U211 ( .B1(n645), .B2(n795), .A(n90), .ZN(n91) );
  AOI21_X1 U212 ( .B1(n789), .B2(n703), .A(n91), .ZN(n801) );
  AOI22_X1 U213 ( .A1(n810), .A2(n266), .B1(n740), .B2(n801), .ZN(n92) );
  OAI211_X1 U214 ( .C1(n833), .C2(n743), .A(n93), .B(n92), .ZN(n94) );
  AOI211_X1 U215 ( .C1(n802), .C2(n774), .A(n95), .B(n94), .ZN(n96) );
  OAI211_X1 U216 ( .C1(n818), .C2(n271), .A(n97), .B(n96), .ZN(data_out[0]) );
  AND2_X1 U217 ( .A1(n607), .A2(data_in[6]), .ZN(n477) );
  AOI21_X1 U218 ( .B1(data_in[13]), .B2(n533), .A(n477), .ZN(n791) );
  NAND2_X1 U219 ( .A1(n607), .A2(data_in[10]), .ZN(n225) );
  NAND2_X1 U220 ( .A1(n729), .A2(n225), .ZN(n108) );
  NAND2_X1 U221 ( .A1(n70), .A2(n108), .ZN(n165) );
  OAI21_X1 U222 ( .B1(n791), .B2(n70), .A(n165), .ZN(n139) );
  INV_X1 U223 ( .A(n139), .ZN(n137) );
  AOI22_X1 U224 ( .A1(n533), .A2(data_in[15]), .B1(n607), .B2(data_in[8]), 
        .ZN(n788) );
  NOR2_X1 U225 ( .A1(n67), .A2(n788), .ZN(n126) );
  AOI22_X1 U226 ( .A1(n533), .A2(data_in[11]), .B1(n607), .B2(data_in[4]), 
        .ZN(n790) );
  NOR2_X1 U227 ( .A1(n790), .A2(n69), .ZN(n676) );
  OAI21_X1 U228 ( .B1(n126), .B2(n676), .A(n62), .ZN(n98) );
  OAI21_X1 U229 ( .B1(n62), .B2(n137), .A(n98), .ZN(n114) );
  AOI22_X1 U230 ( .A1(n533), .A2(data_in[12]), .B1(n607), .B2(data_in[5]), 
        .ZN(n711) );
  INV_X1 U231 ( .A(n711), .ZN(n762) );
  AOI21_X1 U232 ( .B1(n607), .B2(data_in[9]), .A(n99), .ZN(n148) );
  NOR2_X1 U233 ( .A1(n67), .A2(n148), .ZN(n140) );
  AOI21_X1 U234 ( .B1(n63), .B2(n762), .A(n140), .ZN(n135) );
  INV_X1 U235 ( .A(data_in[14]), .ZN(n324) );
  NAND2_X1 U236 ( .A1(n607), .A2(data_in[7]), .ZN(n343) );
  OAI21_X1 U237 ( .B1(n264), .B2(n324), .A(n343), .ZN(n759) );
  INV_X1 U238 ( .A(n759), .ZN(n106) );
  AOI22_X1 U239 ( .A1(n533), .A2(data_in[10]), .B1(n607), .B2(data_in[3]), 
        .ZN(n107) );
  AOI222_X1 U240 ( .A1(n72), .A2(n135), .B1(n106), .B2(n792), .C1(n786), .C2(
        n107), .ZN(n809) );
  NAND2_X1 U241 ( .A1(shift[0]), .A2(n265), .ZN(n814) );
  INV_X1 U242 ( .A(n814), .ZN(n778) );
  NAND2_X1 U243 ( .A1(n70), .A2(n607), .ZN(n340) );
  NOR2_X1 U244 ( .A1(n67), .A2(n104), .ZN(n732) );
  AOI21_X1 U245 ( .B1(data_in[2]), .B2(n333), .A(n732), .ZN(n169) );
  NOR3_X1 U246 ( .A1(n66), .A2(n100), .A3(shift[4]), .ZN(n111) );
  NOR2_X1 U247 ( .A1(n169), .A2(n297), .ZN(n143) );
  NOR2_X1 U248 ( .A1(n64), .A2(n757), .ZN(n307) );
  OAI22_X1 U249 ( .A1(n147), .A2(n795), .B1(n645), .B2(n758), .ZN(n102) );
  AOI211_X1 U250 ( .C1(n789), .C2(n349), .A(n307), .B(n102), .ZN(n822) );
  INV_X1 U251 ( .A(n331), .ZN(n158) );
  OAI22_X1 U252 ( .A1(n365), .A2(n760), .B1(n158), .B2(n795), .ZN(n103) );
  AOI211_X1 U253 ( .C1(n787), .C2(n124), .A(n307), .B(n103), .ZN(n658) );
  NAND2_X1 U254 ( .A1(shift[0]), .A2(n111), .ZN(n827) );
  INV_X1 U255 ( .A(n827), .ZN(n563) );
  NOR2_X1 U256 ( .A1(n67), .A2(n702), .ZN(n302) );
  AOI21_X1 U257 ( .B1(data_in[1]), .B2(n333), .A(n302), .ZN(n142) );
  NOR2_X1 U258 ( .A1(n142), .A2(n792), .ZN(n808) );
  NAND2_X1 U259 ( .A1(n63), .A2(n607), .ZN(n348) );
  NOR2_X1 U260 ( .A1(n69), .A2(n104), .ZN(n541) );
  AOI21_X1 U261 ( .B1(n366), .B2(data_in[2]), .A(n541), .ZN(n163) );
  NOR2_X1 U262 ( .A1(n727), .A2(n63), .ZN(n542) );
  INV_X1 U263 ( .A(n542), .ZN(n105) );
  AOI21_X1 U264 ( .B1(n163), .B2(n105), .A(n534), .ZN(n153) );
  INV_X1 U265 ( .A(n784), .ZN(n812) );
  AOI22_X1 U266 ( .A1(n68), .A2(n148), .B1(n711), .B2(n69), .ZN(n132) );
  NOR2_X1 U267 ( .A1(n106), .A2(n69), .ZN(n121) );
  INV_X1 U268 ( .A(n107), .ZN(n761) );
  NAND2_X1 U269 ( .A1(n69), .A2(n761), .ZN(n696) );
  NAND2_X1 U270 ( .A1(n63), .A2(n108), .ZN(n159) );
  OAI21_X1 U271 ( .B1(n63), .B2(n791), .A(n159), .ZN(n138) );
  NOR2_X1 U272 ( .A1(n788), .A2(n69), .ZN(n129) );
  NOR2_X1 U273 ( .A1(n67), .A2(n790), .ZN(n673) );
  INV_X1 U274 ( .A(n796), .ZN(n112) );
  NAND2_X1 U275 ( .A1(n111), .A2(n258), .ZN(n625) );
  NOR2_X1 U276 ( .A1(n69), .A2(n702), .ZN(n310) );
  AOI21_X1 U277 ( .B1(data_in[1]), .B2(n366), .A(n310), .ZN(n152) );
  OAI21_X1 U278 ( .B1(n699), .B2(n63), .A(n152), .ZN(n117) );
  INV_X1 U279 ( .A(n117), .ZN(n134) );
  AOI221_X1 U280 ( .B1(n705), .B2(n63), .C1(n109), .C2(n69), .A(n62), .ZN(n263) );
  AOI21_X1 U281 ( .B1(n134), .B2(n62), .A(n263), .ZN(n815) );
  INV_X1 U282 ( .A(n637), .ZN(n821) );
  NAND2_X1 U283 ( .A1(n72), .A2(shift[0]), .ZN(n669) );
  NAND2_X1 U284 ( .A1(n553), .A2(n537), .ZN(n545) );
  INV_X1 U285 ( .A(n545), .ZN(n118) );
  NOR2_X1 U286 ( .A1(n605), .A2(n110), .ZN(n800) );
  INV_X1 U287 ( .A(n800), .ZN(n824) );
  NAND2_X1 U288 ( .A1(n111), .A2(n295), .ZN(n136) );
  NAND2_X1 U289 ( .A1(n792), .A2(n349), .ZN(n113) );
  NAND2_X1 U290 ( .A1(n63), .A2(n605), .ZN(n247) );
  OAI211_X1 U291 ( .C1(n147), .C2(n758), .A(n113), .B(n247), .ZN(n683) );
  AOI22_X1 U292 ( .A1(n68), .A2(n645), .B1(data_in[3]), .B2(n366), .ZN(n174)
         );
  NOR2_X1 U293 ( .A1(n69), .A2(n120), .ZN(n649) );
  AOI21_X1 U294 ( .B1(n366), .B2(data_in[11]), .A(n649), .ZN(n171) );
  AOI22_X1 U295 ( .A1(n537), .A2(n705), .B1(n536), .B2(n759), .ZN(n115) );
  OAI222_X1 U296 ( .A1(n534), .A2(n174), .B1(n535), .B2(n171), .C1(n115), .C2(
        n67), .ZN(n164) );
  AOI22_X1 U297 ( .A1(data_in[3]), .A2(n333), .B1(n645), .B2(n69), .ZN(n182)
         );
  INV_X1 U298 ( .A(data_in[11]), .ZN(n119) );
  OAI22_X1 U299 ( .A1(n63), .A2(n120), .B1(n119), .B2(n340), .ZN(n180) );
  OAI21_X1 U300 ( .B1(n121), .B2(n180), .A(n265), .ZN(n122) );
  OAI21_X1 U301 ( .B1(n182), .B2(n297), .A(n122), .ZN(n170) );
  INV_X1 U302 ( .A(n551), .ZN(n715) );
  NAND2_X1 U303 ( .A1(n265), .A2(n258), .ZN(n628) );
  NAND2_X1 U304 ( .A1(n553), .A2(n536), .ZN(n547) );
  INV_X1 U305 ( .A(n547), .ZN(n502) );
  NOR2_X1 U306 ( .A1(n69), .A2(n124), .ZN(n276) );
  AOI21_X1 U307 ( .B1(n681), .B2(data_in[23]), .A(n276), .ZN(n734) );
  INV_X1 U308 ( .A(data_in[19]), .ZN(n455) );
  NOR3_X1 U309 ( .A1(n69), .A2(n264), .A3(n455), .ZN(n680) );
  AOI21_X1 U310 ( .B1(n366), .B2(data_in[12]), .A(n680), .ZN(n125) );
  INV_X1 U311 ( .A(n125), .ZN(n189) );
  OAI21_X1 U312 ( .B1(n126), .B2(n189), .A(n536), .ZN(n127) );
  OAI21_X1 U313 ( .B1(n734), .B2(n534), .A(n127), .ZN(n175) );
  AOI22_X1 U314 ( .A1(n68), .A2(n320), .B1(n333), .B2(data_in[4]), .ZN(n131)
         );
  OAI21_X1 U315 ( .B1(n268), .B2(n340), .A(n128), .ZN(n198) );
  OAI21_X1 U316 ( .B1(n129), .B2(n198), .A(n265), .ZN(n130) );
  OAI21_X1 U317 ( .B1(n131), .B2(n297), .A(n130), .ZN(n183) );
  INV_X1 U318 ( .A(n660), .ZN(n568) );
  AOI22_X1 U319 ( .A1(n792), .A2(n188), .B1(n787), .B2(n331), .ZN(n133) );
  NAND2_X1 U320 ( .A1(n133), .A2(n247), .ZN(n708) );
  NAND2_X1 U321 ( .A1(n265), .A2(n295), .ZN(n651) );
  NOR2_X1 U322 ( .A1(n64), .A2(n787), .ZN(n201) );
  AOI21_X1 U323 ( .B1(n787), .B2(n349), .A(n201), .ZN(n741) );
  INV_X1 U324 ( .A(n651), .ZN(n451) );
  AOI22_X1 U325 ( .A1(n451), .A2(n139), .B1(n568), .B2(n138), .ZN(n145) );
  AOI22_X1 U326 ( .A1(n68), .A2(n147), .B1(n366), .B2(data_in[5]), .ZN(n209)
         );
  AOI21_X1 U327 ( .B1(n607), .B2(data_in[13]), .A(n646), .ZN(n149) );
  NOR2_X1 U328 ( .A1(n149), .A2(n69), .ZN(n207) );
  OAI21_X1 U329 ( .B1(n140), .B2(n207), .A(n536), .ZN(n141) );
  OAI221_X1 U330 ( .B1(n534), .B2(n142), .C1(n534), .C2(n209), .A(n141), .ZN(
        n194) );
  OAI21_X1 U331 ( .B1(n143), .B2(n194), .A(n295), .ZN(n144) );
  OAI211_X1 U332 ( .C1(n834), .C2(n708), .A(n145), .B(n144), .ZN(n146) );
  AOI211_X1 U333 ( .C1(n823), .C2(n741), .A(n800), .B(n146), .ZN(n157) );
  OAI21_X1 U334 ( .B1(n183), .B2(n164), .A(n553), .ZN(n156) );
  OAI21_X1 U335 ( .B1(n175), .B2(n170), .A(n258), .ZN(n155) );
  AOI22_X1 U336 ( .A1(data_in[5]), .A2(n333), .B1(n147), .B2(n69), .ZN(n215)
         );
  NOR2_X1 U337 ( .A1(n148), .A2(n69), .ZN(n150) );
  NOR2_X1 U338 ( .A1(n67), .A2(n149), .ZN(n214) );
  OAI21_X1 U339 ( .B1(n150), .B2(n214), .A(n265), .ZN(n151) );
  OAI221_X1 U340 ( .B1(n297), .B2(n152), .C1(n297), .C2(n215), .A(n151), .ZN(
        n200) );
  OAI21_X1 U341 ( .B1(n153), .B2(n200), .A(n551), .ZN(n154) );
  NAND4_X1 U342 ( .A1(n157), .A2(n156), .A3(n155), .A4(n154), .ZN(data_out[13]) );
  OR2_X1 U343 ( .A1(n188), .A2(n201), .ZN(n768) );
  AOI22_X1 U344 ( .A1(data_in[6]), .A2(n333), .B1(n158), .B2(n69), .ZN(n236)
         );
  INV_X1 U345 ( .A(n159), .ZN(n161) );
  INV_X1 U346 ( .A(n727), .ZN(n160) );
  AOI21_X1 U347 ( .B1(data_in[14]), .B2(n607), .A(n160), .ZN(n166) );
  NOR2_X1 U348 ( .A1(n67), .A2(n166), .ZN(n235) );
  OAI21_X1 U349 ( .B1(n161), .B2(n235), .A(n265), .ZN(n162) );
  OAI221_X1 U350 ( .B1(n297), .B2(n163), .C1(n297), .C2(n236), .A(n162), .ZN(
        n219) );
  NOR2_X1 U351 ( .A1(n69), .A2(n331), .ZN(n731) );
  AOI21_X1 U352 ( .B1(data_in[6]), .B2(n366), .A(n731), .ZN(n226) );
  INV_X1 U353 ( .A(n165), .ZN(n167) );
  NOR2_X1 U354 ( .A1(n166), .A2(n69), .ZN(n224) );
  OAI21_X1 U355 ( .B1(n167), .B2(n224), .A(n536), .ZN(n168) );
  OAI221_X1 U356 ( .B1(n534), .B2(n169), .C1(n534), .C2(n226), .A(n168), .ZN(
        n213) );
  INV_X1 U357 ( .A(n349), .ZN(n178) );
  AOI22_X1 U358 ( .A1(data_in[7]), .A2(n333), .B1(n178), .B2(n69), .ZN(n253)
         );
  AOI21_X1 U359 ( .B1(data_in[15]), .B2(n607), .A(n705), .ZN(n179) );
  NOR2_X1 U360 ( .A1(n67), .A2(n179), .ZN(n251) );
  INV_X1 U361 ( .A(n171), .ZN(n172) );
  OAI21_X1 U362 ( .B1(n251), .B2(n172), .A(n265), .ZN(n173) );
  OAI221_X1 U363 ( .B1(n297), .B2(n174), .C1(n297), .C2(n253), .A(n173), .ZN(
        n240) );
  OAI21_X1 U364 ( .B1(n175), .B2(n240), .A(n551), .ZN(n176) );
  OAI21_X1 U365 ( .B1(n768), .B2(n834), .A(n176), .ZN(n177) );
  AOI211_X1 U366 ( .C1(n64), .C2(n823), .A(n800), .B(n177), .ZN(n187) );
  OAI21_X1 U367 ( .B1(n200), .B2(n213), .A(n258), .ZN(n186) );
  OAI21_X1 U368 ( .B1(n194), .B2(n219), .A(n553), .ZN(n185) );
  AOI22_X1 U369 ( .A1(n68), .A2(n178), .B1(n366), .B2(data_in[7]), .ZN(n252)
         );
  NOR2_X1 U370 ( .A1(n179), .A2(n69), .ZN(n246) );
  OAI21_X1 U371 ( .B1(n246), .B2(n180), .A(n536), .ZN(n181) );
  OAI221_X1 U372 ( .B1(n534), .B2(n182), .C1(n534), .C2(n252), .A(n181), .ZN(
        n234) );
  OAI21_X1 U373 ( .B1(n183), .B2(n234), .A(n295), .ZN(n184) );
  NAND4_X1 U374 ( .A1(n187), .A2(n186), .A3(n185), .A4(n184), .ZN(data_out[15]) );
  OAI21_X1 U375 ( .B1(n375), .B2(n604), .A(n188), .ZN(n196) );
  AND2_X1 U376 ( .A1(n70), .A2(n196), .ZN(n279) );
  AOI21_X1 U377 ( .B1(n366), .B2(data_in[4]), .A(n279), .ZN(n191) );
  AOI22_X1 U378 ( .A1(n533), .A2(data_in[23]), .B1(n607), .B2(data_in[16]), 
        .ZN(n197) );
  NOR2_X1 U379 ( .A1(n67), .A2(n197), .ZN(n275) );
  OAI21_X1 U380 ( .B1(n275), .B2(n189), .A(n265), .ZN(n190) );
  OAI21_X1 U381 ( .B1(n191), .B2(n297), .A(n190), .ZN(n254) );
  NOR3_X1 U382 ( .A1(shift[3]), .A2(n66), .A3(n192), .ZN(n202) );
  NAND2_X1 U383 ( .A1(n202), .A2(n400), .ZN(n481) );
  NOR2_X1 U384 ( .A1(n283), .A2(n201), .ZN(n401) );
  INV_X1 U385 ( .A(n401), .ZN(n364) );
  NAND2_X1 U386 ( .A1(n195), .A2(n69), .ZN(n280) );
  NAND2_X1 U387 ( .A1(n63), .A2(n196), .ZN(n284) );
  NOR2_X1 U388 ( .A1(n197), .A2(n69), .ZN(n281) );
  OAI21_X1 U389 ( .B1(n281), .B2(n198), .A(n536), .ZN(n199) );
  OAI221_X1 U390 ( .B1(n534), .B2(n280), .C1(n534), .C2(n284), .A(n199), .ZN(
        n250) );
  NAND2_X1 U391 ( .A1(n607), .A2(data_in[1]), .ZN(n304) );
  NOR2_X1 U392 ( .A1(n201), .A2(n304), .ZN(n419) );
  NAND2_X1 U393 ( .A1(shift[0]), .A2(n202), .ZN(n523) );
  NAND2_X1 U394 ( .A1(n203), .A2(n64), .ZN(n205) );
  OAI21_X1 U395 ( .B1(n240), .B2(n250), .A(n258), .ZN(n204) );
  OAI211_X1 U396 ( .C1(n364), .C2(n523), .A(n205), .B(n204), .ZN(n206) );
  AOI21_X1 U397 ( .B1(n634), .B2(n419), .A(n206), .ZN(n223) );
  AOI211_X1 U398 ( .C1(n333), .C2(data_in[17]), .A(n302), .B(n207), .ZN(n212)
         );
  INV_X1 U399 ( .A(n265), .ZN(n550) );
  NAND2_X1 U400 ( .A1(n607), .A2(data_in[9]), .ZN(n208) );
  NAND2_X1 U401 ( .A1(n208), .A2(n605), .ZN(n390) );
  INV_X1 U402 ( .A(n390), .ZN(n298) );
  OAI21_X1 U403 ( .B1(n63), .B2(n298), .A(n209), .ZN(n210) );
  INV_X1 U404 ( .A(n210), .ZN(n211) );
  OAI22_X1 U405 ( .A1(n212), .A2(n550), .B1(n211), .B2(n297), .ZN(n278) );
  OAI21_X1 U406 ( .B1(n213), .B2(n278), .A(n551), .ZN(n222) );
  OAI21_X1 U407 ( .B1(n234), .B2(n254), .A(n553), .ZN(n221) );
  AOI211_X1 U408 ( .C1(n366), .C2(data_in[17]), .A(n310), .B(n214), .ZN(n218)
         );
  OAI21_X1 U409 ( .B1(n69), .B2(n298), .A(n215), .ZN(n216) );
  INV_X1 U410 ( .A(n216), .ZN(n217) );
  OAI22_X1 U411 ( .A1(n218), .A2(n535), .B1(n217), .B2(n534), .ZN(n273) );
  OAI21_X1 U412 ( .B1(n219), .B2(n273), .A(n295), .ZN(n220) );
  NAND4_X1 U413 ( .A1(n223), .A2(n222), .A3(n221), .A4(n220), .ZN(data_out[17]) );
  AOI211_X1 U414 ( .C1(data_in[18]), .C2(n333), .A(n732), .B(n224), .ZN(n229)
         );
  NAND2_X1 U415 ( .A1(n605), .A2(n225), .ZN(n571) );
  INV_X1 U416 ( .A(n571), .ZN(n474) );
  OAI21_X1 U417 ( .B1(n63), .B2(n474), .A(n226), .ZN(n227) );
  INV_X1 U418 ( .A(n227), .ZN(n228) );
  OAI22_X1 U419 ( .A1(n229), .A2(n550), .B1(n228), .B2(n297), .ZN(n294) );
  AND2_X1 U420 ( .A1(n607), .A2(data_in[2]), .ZN(n532) );
  NOR2_X1 U421 ( .A1(n64), .A2(n532), .ZN(n231) );
  INV_X1 U422 ( .A(n231), .ZN(n442) );
  AOI21_X1 U423 ( .B1(n823), .B2(n442), .A(n800), .ZN(n334) );
  OAI21_X1 U424 ( .B1(n320), .B2(n795), .A(n247), .ZN(n230) );
  AOI21_X1 U425 ( .B1(n787), .B2(n231), .A(n230), .ZN(n443) );
  AOI22_X1 U426 ( .A1(n634), .A2(n443), .B1(n632), .B2(n419), .ZN(n232) );
  OAI211_X1 U427 ( .C1(n834), .C2(n605), .A(n334), .B(n232), .ZN(n233) );
  AOI221_X1 U428 ( .B1(n234), .B2(n551), .C1(n294), .C2(n551), .A(n233), .ZN(
        n244) );
  OAI21_X1 U429 ( .B1(n254), .B2(n273), .A(n258), .ZN(n243) );
  OAI21_X1 U430 ( .B1(n250), .B2(n278), .A(n553), .ZN(n242) );
  AOI211_X1 U431 ( .C1(data_in[18]), .C2(n366), .A(n541), .B(n235), .ZN(n239)
         );
  OAI21_X1 U432 ( .B1(n69), .B2(n474), .A(n236), .ZN(n237) );
  INV_X1 U433 ( .A(n237), .ZN(n238) );
  OAI22_X1 U434 ( .A1(n239), .A2(n535), .B1(n238), .B2(n534), .ZN(n296) );
  OAI21_X1 U435 ( .B1(n240), .B2(n296), .A(n295), .ZN(n241) );
  NAND4_X1 U436 ( .A1(n244), .A2(n243), .A3(n242), .A4(n241), .ZN(data_out[18]) );
  AOI21_X1 U437 ( .B1(data_in[3]), .B2(n607), .A(n64), .ZN(n441) );
  AOI21_X1 U438 ( .B1(n802), .B2(n442), .A(n800), .ZN(n245) );
  OAI21_X1 U439 ( .B1(n441), .B2(n668), .A(n245), .ZN(n356) );
  OAI22_X1 U440 ( .A1(n63), .A2(n707), .B1(n340), .B2(n455), .ZN(n350) );
  NOR2_X1 U441 ( .A1(n246), .A2(n350), .ZN(n328) );
  NOR2_X1 U442 ( .A1(n550), .A2(n715), .ZN(n623) );
  INV_X1 U443 ( .A(n623), .ZN(n678) );
  AOI22_X1 U444 ( .A1(n792), .A2(n304), .B1(n787), .B2(n441), .ZN(n248) );
  NAND2_X1 U445 ( .A1(n248), .A2(n247), .ZN(n472) );
  OAI22_X1 U446 ( .A1(n328), .A2(n678), .B1(n481), .B2(n472), .ZN(n249) );
  AOI211_X1 U447 ( .C1(n551), .C2(n250), .A(n356), .B(n249), .ZN(n261) );
  OAI22_X1 U448 ( .A1(n69), .A2(n707), .B1(n455), .B2(n348), .ZN(n341) );
  NOR2_X1 U449 ( .A1(n251), .A2(n341), .ZN(n327) );
  INV_X1 U450 ( .A(n295), .ZN(n718) );
  NOR2_X1 U451 ( .A1(n535), .A2(n718), .ZN(n514) );
  INV_X1 U452 ( .A(n514), .ZN(n677) );
  NOR2_X1 U453 ( .A1(n297), .A2(n715), .ZN(n621) );
  AOI21_X1 U454 ( .B1(data_in[11]), .B2(n607), .A(n64), .ZN(n629) );
  OAI21_X1 U455 ( .B1(n63), .B2(n629), .A(n252), .ZN(n299) );
  AOI22_X1 U456 ( .A1(n632), .A2(n443), .B1(n621), .B2(n299), .ZN(n256) );
  NAND2_X1 U457 ( .A1(n537), .A2(n295), .ZN(n650) );
  INV_X1 U458 ( .A(n650), .ZN(n682) );
  OAI21_X1 U459 ( .B1(n629), .B2(n70), .A(n253), .ZN(n301) );
  AOI22_X1 U460 ( .A1(n295), .A2(n254), .B1(n682), .B2(n301), .ZN(n255) );
  OAI211_X1 U461 ( .C1(n327), .C2(n677), .A(n256), .B(n255), .ZN(n257) );
  AOI221_X1 U462 ( .B1(n273), .B2(n553), .C1(n294), .C2(n553), .A(n257), .ZN(
        n260) );
  OAI21_X1 U463 ( .B1(n278), .B2(n296), .A(n258), .ZN(n259) );
  NAND3_X1 U464 ( .A1(n261), .A2(n260), .A3(n259), .ZN(data_out[19]) );
  AOI211_X1 U465 ( .C1(n646), .C2(n69), .A(n310), .B(n72), .ZN(n262) );
  NOR2_X1 U466 ( .A1(n263), .A2(n262), .ZN(n544) );
  OAI21_X1 U467 ( .B1(n375), .B2(n264), .A(n304), .ZN(n756) );
  NAND3_X1 U468 ( .A1(n70), .A2(n756), .A3(n265), .ZN(n691) );
  INV_X1 U469 ( .A(n691), .ZN(n552) );
  INV_X1 U470 ( .A(n756), .ZN(n713) );
  OAI22_X1 U471 ( .A1(n713), .A2(n535), .B1(n534), .B2(n697), .ZN(n270) );
  OAI22_X1 U472 ( .A1(n268), .A2(n534), .B1(n267), .B2(n535), .ZN(n269) );
  AOI22_X1 U473 ( .A1(n68), .A2(n270), .B1(n681), .B2(n269), .ZN(n670) );
  AOI22_X1 U474 ( .A1(n553), .A2(n296), .B1(n551), .B2(n273), .ZN(n293) );
  AOI21_X1 U475 ( .B1(data_in[4]), .B2(n607), .A(n64), .ZN(n491) );
  INV_X1 U476 ( .A(n491), .ZN(n512) );
  AOI21_X1 U477 ( .B1(n823), .B2(n512), .A(n800), .ZN(n274) );
  OAI21_X1 U478 ( .B1(n441), .B2(n834), .A(n274), .ZN(n369) );
  NOR2_X1 U479 ( .A1(n276), .A2(n275), .ZN(n323) );
  OAI22_X1 U480 ( .A1(n323), .A2(n677), .B1(n523), .B2(n472), .ZN(n277) );
  AOI211_X1 U481 ( .C1(n295), .C2(n278), .A(n369), .B(n277), .ZN(n292) );
  NOR2_X1 U482 ( .A1(n669), .A2(n550), .ZN(n593) );
  INV_X1 U483 ( .A(n593), .ZN(n709) );
  OAI22_X1 U484 ( .A1(n327), .A2(n719), .B1(n328), .B2(n709), .ZN(n290) );
  AOI21_X1 U485 ( .B1(n607), .B2(data_in[12]), .A(n64), .ZN(n473) );
  INV_X1 U486 ( .A(n473), .ZN(n570) );
  NOR2_X1 U487 ( .A1(n279), .A2(n570), .ZN(n329) );
  INV_X1 U488 ( .A(data_in[20]), .ZN(n484) );
  OAI21_X1 U489 ( .B1(n484), .B2(n340), .A(n280), .ZN(n372) );
  NOR2_X1 U490 ( .A1(n281), .A2(n372), .ZN(n363) );
  OAI22_X1 U491 ( .A1(n329), .A2(n650), .B1(n363), .B2(n678), .ZN(n289) );
  INV_X1 U492 ( .A(n294), .ZN(n287) );
  OAI22_X1 U493 ( .A1(n795), .A2(n442), .B1(n758), .B2(n512), .ZN(n282) );
  AOI211_X1 U494 ( .C1(n789), .C2(n283), .A(n307), .B(n282), .ZN(n511) );
  OAI21_X1 U495 ( .B1(n63), .B2(n473), .A(n284), .ZN(n325) );
  AOI22_X1 U496 ( .A1(n634), .A2(n511), .B1(n621), .B2(n325), .ZN(n286) );
  NOR2_X1 U497 ( .A1(n669), .A2(n297), .ZN(n303) );
  INV_X1 U498 ( .A(n684), .ZN(n701) );
  AOI22_X1 U499 ( .A1(n303), .A2(n299), .B1(n701), .B2(n301), .ZN(n285) );
  OAI211_X1 U500 ( .C1(n287), .C2(n671), .A(n286), .B(n285), .ZN(n288) );
  NOR3_X1 U501 ( .A1(n290), .A2(n289), .A3(n288), .ZN(n291) );
  NAND3_X1 U502 ( .A1(n293), .A2(n292), .A3(n291), .ZN(data_out[20]) );
  AOI22_X1 U503 ( .A1(n551), .A2(n296), .B1(n295), .B2(n294), .ZN(n319) );
  NOR2_X1 U504 ( .A1(n297), .A2(shift[0]), .ZN(n807) );
  INV_X1 U505 ( .A(n807), .ZN(n797) );
  AOI21_X1 U506 ( .B1(data_in[13]), .B2(n607), .A(n64), .ZN(n395) );
  AOI22_X1 U507 ( .A1(n787), .A2(n395), .B1(n298), .B2(n789), .ZN(n509) );
  OAI21_X1 U508 ( .B1(n71), .B2(n299), .A(n509), .ZN(n326) );
  INV_X1 U509 ( .A(n776), .ZN(n816) );
  NOR2_X1 U510 ( .A1(n795), .A2(n390), .ZN(n453) );
  INV_X1 U511 ( .A(n453), .ZN(n300) );
  NAND2_X1 U512 ( .A1(n786), .A2(n395), .ZN(n458) );
  OAI211_X1 U513 ( .C1(n62), .C2(n301), .A(n300), .B(n458), .ZN(n337) );
  OAI22_X1 U514 ( .A1(n797), .A2(n326), .B1(n816), .B2(n337), .ZN(n317) );
  OAI22_X1 U515 ( .A1(n327), .A2(n547), .B1(n323), .B2(n719), .ZN(n316) );
  OAI22_X1 U516 ( .A1(n328), .A2(n628), .B1(n363), .B2(n709), .ZN(n315) );
  INV_X1 U517 ( .A(data_in[21]), .ZN(n309) );
  OAI22_X1 U518 ( .A1(n69), .A2(n703), .B1(n348), .B2(n309), .ZN(n405) );
  AOI211_X1 U519 ( .C1(n333), .C2(data_in[17]), .A(n302), .B(n405), .ZN(n378)
         );
  AOI22_X1 U520 ( .A1(n632), .A2(n511), .B1(n303), .B2(n325), .ZN(n313) );
  INV_X1 U521 ( .A(n304), .ZN(n344) );
  OAI21_X1 U522 ( .B1(n305), .B2(n604), .A(n605), .ZN(n586) );
  OAI22_X1 U523 ( .A1(n344), .A2(n760), .B1(n758), .B2(n586), .ZN(n306) );
  AOI211_X1 U524 ( .C1(n792), .C2(n441), .A(n307), .B(n306), .ZN(n564) );
  AOI22_X1 U525 ( .A1(n802), .A2(n512), .B1(n823), .B2(n586), .ZN(n308) );
  NAND2_X1 U526 ( .A1(n308), .A2(n824), .ZN(n389) );
  OAI22_X1 U527 ( .A1(n63), .A2(n703), .B1(n309), .B2(n340), .ZN(n396) );
  AOI211_X1 U528 ( .C1(n366), .C2(data_in[17]), .A(n310), .B(n396), .ZN(n379)
         );
  OAI22_X1 U529 ( .A1(n329), .A2(n684), .B1(n379), .B2(n678), .ZN(n311) );
  AOI211_X1 U530 ( .C1(n634), .C2(n564), .A(n389), .B(n311), .ZN(n312) );
  OAI211_X1 U531 ( .C1(n378), .C2(n677), .A(n313), .B(n312), .ZN(n314) );
  NOR4_X1 U532 ( .A1(n317), .A2(n316), .A3(n315), .A4(n314), .ZN(n318) );
  NAND2_X1 U533 ( .A1(n319), .A2(n318), .ZN(data_out[21]) );
  AOI22_X1 U534 ( .A1(n320), .A2(n786), .B1(n787), .B2(n477), .ZN(n322) );
  AOI22_X1 U535 ( .A1(n792), .A2(n512), .B1(n789), .B2(n442), .ZN(n321) );
  NAND2_X1 U536 ( .A1(n322), .A2(n321), .ZN(n618) );
  INV_X1 U537 ( .A(n323), .ZN(n339) );
  OAI21_X1 U538 ( .B1(n324), .B2(n604), .A(n605), .ZN(n569) );
  OAI222_X1 U539 ( .A1(n760), .A2(n571), .B1(n325), .B2(n72), .C1(n758), .C2(
        n569), .ZN(n354) );
  AOI21_X1 U540 ( .B1(n474), .B2(n792), .A(n329), .ZN(n330) );
  INV_X1 U541 ( .A(n330), .ZN(n342) );
  OAI22_X1 U542 ( .A1(n63), .A2(n331), .B1(n576), .B2(n340), .ZN(n421) );
  AOI211_X1 U543 ( .C1(data_in[18]), .C2(n366), .A(n541), .B(n421), .ZN(n403)
         );
  OAI22_X1 U544 ( .A1(n363), .A2(n628), .B1(n403), .B2(n678), .ZN(n336) );
  AOI21_X1 U545 ( .B1(data_in[22]), .B2(n366), .A(n731), .ZN(n332) );
  INV_X1 U546 ( .A(n332), .ZN(n416) );
  AOI211_X1 U547 ( .C1(data_in[18]), .C2(n333), .A(n732), .B(n416), .ZN(n406)
         );
  NAND2_X1 U548 ( .A1(n802), .A2(n586), .ZN(n415) );
  OAI211_X1 U549 ( .C1(n406), .C2(n677), .A(n334), .B(n415), .ZN(n335) );
  OAI22_X1 U550 ( .A1(n403), .A2(n709), .B1(n406), .B2(n719), .ZN(n338) );
  AOI21_X1 U551 ( .B1(n568), .B2(n339), .A(n338), .ZN(n362) );
  OAI22_X1 U552 ( .A1(n68), .A2(n349), .B1(n347), .B2(n340), .ZN(n446) );
  NOR2_X1 U553 ( .A1(n341), .A2(n446), .ZN(n404) );
  INV_X1 U554 ( .A(n404), .ZN(n423) );
  OAI22_X1 U555 ( .A1(n379), .A2(n628), .B1(n637), .B2(n342), .ZN(n360) );
  NAND2_X1 U556 ( .A1(n343), .A2(n605), .ZN(n587) );
  OAI22_X1 U557 ( .A1(n344), .A2(n757), .B1(n758), .B2(n587), .ZN(n345) );
  AOI21_X1 U558 ( .B1(n789), .B2(n441), .A(n345), .ZN(n346) );
  OAI21_X1 U559 ( .B1(n795), .B2(n586), .A(n346), .ZN(n615) );
  OAI22_X1 U560 ( .A1(n69), .A2(n349), .B1(n348), .B2(n347), .ZN(n445) );
  NOR2_X1 U561 ( .A1(n350), .A2(n445), .ZN(n428) );
  OAI22_X1 U562 ( .A1(n378), .A2(n547), .B1(n428), .B2(n677), .ZN(n351) );
  AOI21_X1 U563 ( .B1(n632), .B2(n618), .A(n351), .ZN(n358) );
  AOI21_X1 U564 ( .B1(data_in[15]), .B2(n607), .A(n64), .ZN(n585) );
  AOI22_X1 U565 ( .A1(n792), .A2(n395), .B1(n787), .B2(n585), .ZN(n352) );
  OAI21_X1 U566 ( .B1(n390), .B2(n757), .A(n352), .ZN(n353) );
  AOI21_X1 U567 ( .B1(n789), .B2(n629), .A(n353), .ZN(n633) );
  OAI22_X1 U568 ( .A1(n629), .A2(n816), .B1(n827), .B2(n354), .ZN(n355) );
  AOI211_X1 U569 ( .C1(n633), .C2(n807), .A(n356), .B(n355), .ZN(n357) );
  OAI211_X1 U570 ( .C1(n481), .C2(n615), .A(n358), .B(n357), .ZN(n359) );
  AOI211_X1 U571 ( .C1(n623), .C2(n423), .A(n360), .B(n359), .ZN(n361) );
  OAI211_X1 U572 ( .C1(n363), .C2(n651), .A(n362), .B(n361), .ZN(data_out[23])
         );
  AOI21_X1 U573 ( .B1(data_in[16]), .B2(n607), .A(n64), .ZN(n638) );
  NOR2_X1 U574 ( .A1(n638), .A2(n816), .ZN(n581) );
  NAND3_X1 U575 ( .A1(shift[3]), .A2(shift_type[0]), .A3(shift[4]), .ZN(n399)
         );
  NOR2_X1 U576 ( .A1(shift[0]), .A2(n399), .ZN(n566) );
  INV_X1 U577 ( .A(n566), .ZN(n614) );
  OAI22_X1 U578 ( .A1(n629), .A2(n637), .B1(n364), .B2(n614), .ZN(n368) );
  AOI21_X1 U579 ( .B1(data_in[24]), .B2(n607), .A(n365), .ZN(n470) );
  NOR2_X1 U580 ( .A1(n67), .A2(n470), .ZN(n492) );
  AOI21_X1 U581 ( .B1(data_in[20]), .B2(n366), .A(n492), .ZN(n449) );
  OAI22_X1 U582 ( .A1(n403), .A2(n628), .B1(n449), .B2(n678), .ZN(n367) );
  NOR4_X1 U583 ( .A1(n581), .A2(n369), .A3(n368), .A4(n367), .ZN(n386) );
  NOR2_X1 U584 ( .A1(n760), .A2(n570), .ZN(n371) );
  OAI22_X1 U585 ( .A1(n795), .A2(n569), .B1(n571), .B2(n757), .ZN(n370) );
  AOI211_X1 U586 ( .C1(n638), .C2(n787), .A(n371), .B(n370), .ZN(n398) );
  AOI22_X1 U587 ( .A1(n563), .A2(n633), .B1(n807), .B2(n398), .ZN(n385) );
  INV_X1 U588 ( .A(n470), .ZN(n373) );
  AOI21_X1 U589 ( .B1(n373), .B2(n68), .A(n372), .ZN(n444) );
  OAI22_X1 U590 ( .A1(n547), .A2(n406), .B1(n677), .B2(n444), .ZN(n374) );
  INV_X1 U591 ( .A(n374), .ZN(n384) );
  OAI21_X1 U592 ( .B1(n375), .B2(n604), .A(n605), .ZN(n582) );
  INV_X1 U593 ( .A(n582), .ZN(n610) );
  OAI22_X1 U594 ( .A1(n477), .A2(n795), .B1(n442), .B2(n757), .ZN(n376) );
  AOI21_X1 U595 ( .B1(n787), .B2(n610), .A(n376), .ZN(n377) );
  OAI21_X1 U596 ( .B1(n760), .B2(n512), .A(n377), .ZN(n387) );
  OAI22_X1 U597 ( .A1(n481), .A2(n387), .B1(n523), .B2(n615), .ZN(n382) );
  OAI22_X1 U598 ( .A1(n378), .A2(n660), .B1(n428), .B2(n719), .ZN(n381) );
  OAI22_X1 U599 ( .A1(n379), .A2(n651), .B1(n404), .B2(n709), .ZN(n380) );
  NOR3_X1 U600 ( .A1(n382), .A2(n381), .A3(n380), .ZN(n383) );
  NAND4_X1 U601 ( .A1(n386), .A2(n385), .A3(n384), .A4(n383), .ZN(data_out[24]) );
  AOI21_X1 U602 ( .B1(n607), .B2(data_in[17]), .A(n64), .ZN(n456) );
  INV_X1 U603 ( .A(n456), .ZN(n527) );
  OAI22_X1 U604 ( .A1(n638), .A2(n637), .B1(n523), .B2(n387), .ZN(n388) );
  AOI211_X1 U605 ( .C1(n776), .C2(n527), .A(n389), .B(n388), .ZN(n414) );
  NOR2_X1 U606 ( .A1(n760), .A2(n586), .ZN(n392) );
  OAI22_X1 U607 ( .A1(n795), .A2(n587), .B1(n758), .B2(n390), .ZN(n391) );
  AOI211_X1 U608 ( .C1(n441), .C2(n786), .A(n392), .B(n391), .ZN(n438) );
  AOI22_X1 U609 ( .A1(n792), .A2(n585), .B1(n786), .B2(n629), .ZN(n393) );
  OAI21_X1 U610 ( .B1(n758), .B2(n527), .A(n393), .ZN(n394) );
  AOI21_X1 U611 ( .B1(n789), .B2(n395), .A(n394), .ZN(n427) );
  AOI22_X1 U612 ( .A1(n634), .A2(n438), .B1(n807), .B2(n427), .ZN(n413) );
  AOI21_X1 U613 ( .B1(data_in[25]), .B2(n607), .A(n64), .ZN(n596) );
  INV_X1 U614 ( .A(n396), .ZN(n397) );
  OAI21_X1 U615 ( .B1(n596), .B2(n70), .A(n397), .ZN(n497) );
  AOI22_X1 U616 ( .A1(n563), .A2(n398), .B1(n514), .B2(n497), .ZN(n412) );
  NOR2_X1 U617 ( .A1(n400), .A2(n399), .ZN(n619) );
  AOI22_X1 U618 ( .A1(n401), .A2(n619), .B1(n419), .B2(n566), .ZN(n402) );
  OAI21_X1 U619 ( .B1(n403), .B2(n651), .A(n402), .ZN(n410) );
  OAI22_X1 U620 ( .A1(n404), .A2(n628), .B1(n449), .B2(n709), .ZN(n409) );
  OAI22_X1 U621 ( .A1(n428), .A2(n547), .B1(n444), .B2(n719), .ZN(n408) );
  INV_X1 U622 ( .A(n596), .ZN(n513) );
  AOI21_X1 U623 ( .B1(n69), .B2(n513), .A(n405), .ZN(n467) );
  OAI22_X1 U624 ( .A1(n406), .A2(n660), .B1(n467), .B2(n678), .ZN(n407) );
  NOR4_X1 U625 ( .A1(n410), .A2(n409), .A3(n408), .A4(n407), .ZN(n411) );
  NAND4_X1 U626 ( .A1(n414), .A2(n413), .A3(n412), .A4(n411), .ZN(data_out[25]) );
  NAND2_X1 U627 ( .A1(n776), .A2(n569), .ZN(n489) );
  OAI211_X1 U628 ( .C1(n474), .C2(n668), .A(n415), .B(n489), .ZN(n418) );
  AOI21_X1 U629 ( .B1(data_in[26]), .B2(n607), .A(n64), .ZN(n591) );
  INV_X1 U630 ( .A(n591), .ZN(n422) );
  AOI21_X1 U631 ( .B1(n69), .B2(n422), .A(n416), .ZN(n506) );
  OAI22_X1 U632 ( .A1(n467), .A2(n709), .B1(n506), .B2(n678), .ZN(n417) );
  AOI211_X1 U633 ( .C1(n821), .C2(n527), .A(n418), .B(n417), .ZN(n440) );
  INV_X1 U634 ( .A(n740), .ZN(n767) );
  AOI22_X1 U635 ( .A1(n419), .A2(n619), .B1(n443), .B2(n566), .ZN(n420) );
  NAND2_X1 U636 ( .A1(n765), .A2(n442), .ZN(n583) );
  OAI211_X1 U637 ( .C1(n767), .C2(n605), .A(n420), .B(n583), .ZN(n437) );
  AOI21_X1 U638 ( .B1(n422), .B2(n68), .A(n421), .ZN(n466) );
  INV_X1 U639 ( .A(n466), .ZN(n526) );
  AOI22_X1 U640 ( .A1(n451), .A2(n423), .B1(n514), .B2(n526), .ZN(n435) );
  INV_X1 U641 ( .A(n444), .ZN(n424) );
  AOI22_X1 U642 ( .A1(n502), .A2(n424), .B1(n493), .B2(n497), .ZN(n434) );
  NAND2_X1 U643 ( .A1(n607), .A2(data_in[18]), .ZN(n574) );
  AOI22_X1 U644 ( .A1(n787), .A2(n574), .B1(n786), .B2(n473), .ZN(n425) );
  OAI21_X1 U645 ( .B1(n760), .B2(n569), .A(n425), .ZN(n426) );
  AOI21_X1 U646 ( .B1(n792), .B2(n638), .A(n426), .ZN(n460) );
  AOI22_X1 U647 ( .A1(n563), .A2(n427), .B1(n807), .B2(n460), .ZN(n433) );
  INV_X1 U648 ( .A(n428), .ZN(n431) );
  OAI22_X1 U649 ( .A1(n758), .A2(n571), .B1(n757), .B2(n512), .ZN(n430) );
  OAI22_X1 U650 ( .A1(n477), .A2(n760), .B1(n795), .B2(n582), .ZN(n429) );
  NOR2_X1 U651 ( .A1(n430), .A2(n429), .ZN(n454) );
  AOI22_X1 U652 ( .A1(n568), .A2(n431), .B1(n634), .B2(n454), .ZN(n432) );
  NAND4_X1 U653 ( .A1(n435), .A2(n434), .A3(n433), .A4(n432), .ZN(n436) );
  AOI211_X1 U654 ( .C1(n632), .C2(n438), .A(n437), .B(n436), .ZN(n439) );
  OAI211_X1 U655 ( .C1(n449), .C2(n628), .A(n440), .B(n439), .ZN(data_out[26])
         );
  INV_X1 U656 ( .A(n441), .ZN(n488) );
  AOI22_X1 U657 ( .A1(n765), .A2(n488), .B1(n740), .B2(n442), .ZN(n644) );
  NAND2_X1 U658 ( .A1(n821), .A2(n569), .ZN(n504) );
  AOI21_X1 U659 ( .B1(data_in[27]), .B2(n607), .A(n64), .ZN(n448) );
  INV_X1 U660 ( .A(n448), .ZN(n622) );
  AOI21_X1 U661 ( .B1(n69), .B2(n622), .A(n445), .ZN(n579) );
  INV_X1 U662 ( .A(n446), .ZN(n447) );
  OAI21_X1 U663 ( .B1(n448), .B2(n70), .A(n447), .ZN(n567) );
  AOI22_X1 U664 ( .A1(n502), .A2(n497), .B1(n514), .B2(n567), .ZN(n464) );
  INV_X1 U665 ( .A(n449), .ZN(n450) );
  AOI22_X1 U666 ( .A1(n451), .A2(n450), .B1(n493), .B2(n526), .ZN(n463) );
  OAI22_X1 U667 ( .A1(n757), .A2(n586), .B1(n760), .B2(n587), .ZN(n452) );
  AOI211_X1 U668 ( .C1(n629), .C2(n787), .A(n453), .B(n452), .ZN(n479) );
  AOI22_X1 U669 ( .A1(n634), .A2(n479), .B1(n632), .B2(n454), .ZN(n462) );
  NOR2_X1 U670 ( .A1(n455), .A2(n604), .ZN(n620) );
  AOI22_X1 U671 ( .A1(n792), .A2(n456), .B1(n789), .B2(n585), .ZN(n457) );
  OAI211_X1 U672 ( .C1(n758), .C2(n620), .A(n458), .B(n457), .ZN(n459) );
  INV_X1 U673 ( .A(n459), .ZN(n478) );
  AOI22_X1 U674 ( .A1(n563), .A2(n460), .B1(n807), .B2(n478), .ZN(n461) );
  NAND4_X1 U675 ( .A1(n464), .A2(n463), .A3(n462), .A4(n461), .ZN(n465) );
  OAI22_X1 U676 ( .A1(n651), .A2(n467), .B1(n547), .B2(n466), .ZN(n468) );
  INV_X1 U677 ( .A(n468), .ZN(n501) );
  AOI221_X1 U678 ( .B1(n470), .B2(n63), .C1(n469), .C2(n69), .A(n604), .ZN(
        n589) );
  INV_X1 U679 ( .A(n579), .ZN(n471) );
  AOI22_X1 U680 ( .A1(n623), .A2(n589), .B1(n593), .B2(n471), .ZN(n500) );
  INV_X1 U681 ( .A(n619), .ZN(n517) );
  OAI22_X1 U682 ( .A1(n629), .A2(n834), .B1(n472), .B2(n517), .ZN(n483) );
  AOI22_X1 U683 ( .A1(n787), .A2(n473), .B1(n789), .B2(n610), .ZN(n476) );
  NAND2_X1 U684 ( .A1(n792), .A2(n474), .ZN(n475) );
  OAI211_X1 U685 ( .C1(n477), .C2(n757), .A(n476), .B(n475), .ZN(n522) );
  AOI22_X1 U686 ( .A1(n632), .A2(n479), .B1(n563), .B2(n478), .ZN(n480) );
  OAI21_X1 U687 ( .B1(n481), .B2(n522), .A(n480), .ZN(n482) );
  AOI211_X1 U688 ( .C1(n823), .C2(n570), .A(n483), .B(n482), .ZN(n499) );
  NOR2_X1 U689 ( .A1(n585), .A2(n637), .ZN(n487) );
  AOI221_X1 U690 ( .B1(n638), .B2(n63), .C1(n484), .C2(n69), .A(n604), .ZN(
        n578) );
  INV_X1 U691 ( .A(n574), .ZN(n485) );
  OAI222_X1 U692 ( .A1(n757), .A2(n569), .B1(n62), .B2(n578), .C1(n795), .C2(
        n485), .ZN(n531) );
  OAI22_X1 U693 ( .A1(n506), .A2(n628), .B1(n797), .B2(n531), .ZN(n486) );
  AOI211_X1 U694 ( .C1(n740), .C2(n488), .A(n487), .B(n486), .ZN(n490) );
  OAI211_X1 U695 ( .C1(n491), .C2(n743), .A(n490), .B(n489), .ZN(n496) );
  NOR2_X1 U696 ( .A1(n64), .A2(n492), .ZN(n561) );
  AOI22_X1 U697 ( .A1(n493), .A2(n567), .B1(n511), .B2(n566), .ZN(n494) );
  OAI21_X1 U698 ( .B1(n561), .B2(n677), .A(n494), .ZN(n495) );
  AOI211_X1 U699 ( .C1(n568), .C2(n497), .A(n496), .B(n495), .ZN(n498) );
  NAND4_X1 U700 ( .A1(n501), .A2(n500), .A3(n499), .A4(n498), .ZN(data_out[28]) );
  AOI22_X1 U701 ( .A1(n502), .A2(n567), .B1(n564), .B2(n566), .ZN(n503) );
  OAI21_X1 U702 ( .B1(n561), .B2(n719), .A(n503), .ZN(n525) );
  AOI22_X1 U703 ( .A1(n802), .A2(n570), .B1(n765), .B2(n586), .ZN(n505) );
  OAI211_X1 U704 ( .C1(n585), .C2(n816), .A(n505), .B(n504), .ZN(n508) );
  OAI22_X1 U705 ( .A1(n579), .A2(n628), .B1(n506), .B2(n651), .ZN(n507) );
  AOI211_X1 U706 ( .C1(n593), .C2(n589), .A(n508), .B(n507), .ZN(n521) );
  OAI21_X1 U707 ( .B1(n757), .B2(n587), .A(n509), .ZN(n510) );
  AOI21_X1 U708 ( .B1(n792), .B2(n629), .A(n510), .ZN(n565) );
  INV_X1 U709 ( .A(n511), .ZN(n518) );
  AOI22_X1 U710 ( .A1(n823), .A2(n587), .B1(n740), .B2(n512), .ZN(n516) );
  OAI221_X1 U711 ( .B1(n513), .B2(n69), .C1(data_in[29]), .C2(n63), .A(n607), 
        .ZN(n627) );
  INV_X1 U712 ( .A(n627), .ZN(n592) );
  AOI22_X1 U713 ( .A1(n623), .A2(n592), .B1(n514), .B2(n513), .ZN(n515) );
  OAI211_X1 U714 ( .C1(n518), .C2(n517), .A(n516), .B(n515), .ZN(n519) );
  AOI21_X1 U715 ( .B1(n634), .B2(n565), .A(n519), .ZN(n520) );
  OAI211_X1 U716 ( .C1(n523), .C2(n522), .A(n521), .B(n520), .ZN(n524) );
  AOI211_X1 U717 ( .C1(n568), .C2(n526), .A(n525), .B(n524), .ZN(n530) );
  OAI221_X1 U718 ( .B1(n63), .B2(data_in[21]), .C1(n70), .C2(n527), .A(n607), 
        .ZN(n624) );
  INV_X1 U719 ( .A(n620), .ZN(n528) );
  AOI222_X1 U720 ( .A1(n624), .A2(n71), .B1(n585), .B2(n786), .C1(n528), .C2(
        n792), .ZN(n562) );
  NAND2_X1 U721 ( .A1(n807), .A2(n562), .ZN(n529) );
  AOI21_X1 U722 ( .B1(data_in[9]), .B2(n533), .A(n532), .ZN(n785) );
  OAI22_X1 U723 ( .A1(n785), .A2(n535), .B1(n534), .B2(n729), .ZN(n540) );
  AOI22_X1 U724 ( .A1(n537), .A2(data_in[13]), .B1(n536), .B2(data_in[5]), 
        .ZN(n538) );
  INV_X1 U725 ( .A(n538), .ZN(n539) );
  AOI22_X1 U726 ( .A1(n68), .A2(n540), .B1(n681), .B2(n539), .ZN(n716) );
  NOR2_X1 U727 ( .A1(n542), .A2(n541), .ZN(n679) );
  AOI22_X1 U728 ( .A1(n62), .A2(n679), .B1(n543), .B2(n72), .ZN(n656) );
  AOI22_X1 U729 ( .A1(n802), .A2(n544), .B1(n823), .B2(n656), .ZN(n560) );
  OAI22_X1 U730 ( .A1(n653), .A2(n545), .B1(n674), .B2(n628), .ZN(n558) );
  AOI22_X1 U731 ( .A1(n658), .A2(n765), .B1(n822), .B2(n740), .ZN(n546) );
  OAI21_X1 U732 ( .B1(n661), .B2(n547), .A(n546), .ZN(n557) );
  OAI22_X1 U733 ( .A1(n549), .A2(n660), .B1(n548), .B2(n652), .ZN(n556) );
  NOR3_X1 U734 ( .A1(n67), .A2(n785), .A3(n550), .ZN(n657) );
  AOI22_X1 U735 ( .A1(n553), .A2(n552), .B1(n551), .B2(n657), .ZN(n554) );
  OAI21_X1 U736 ( .B1(n670), .B2(n671), .A(n554), .ZN(n555) );
  NOR4_X1 U737 ( .A1(n558), .A2(n557), .A3(n556), .A4(n555), .ZN(n559) );
  OAI211_X1 U738 ( .C1(n716), .C2(n718), .A(n560), .B(n559), .ZN(data_out[2])
         );
  AOI21_X1 U739 ( .B1(n792), .B2(n591), .A(n561), .ZN(n613) );
  AOI22_X1 U740 ( .A1(n782), .A2(n613), .B1(n563), .B2(n562), .ZN(n602) );
  AOI22_X1 U741 ( .A1(n632), .A2(n565), .B1(n564), .B2(n619), .ZN(n601) );
  AOI22_X1 U742 ( .A1(n568), .A2(n567), .B1(n566), .B2(n618), .ZN(n600) );
  AOI22_X1 U743 ( .A1(n792), .A2(n570), .B1(n787), .B2(n569), .ZN(n573) );
  NAND2_X1 U744 ( .A1(n789), .A2(n571), .ZN(n572) );
  OAI211_X1 U745 ( .C1(n610), .C2(n757), .A(n573), .B(n572), .ZN(n631) );
  NOR2_X1 U746 ( .A1(n604), .A2(n758), .ZN(n588) );
  INV_X1 U747 ( .A(n588), .ZN(n575) );
  OAI22_X1 U748 ( .A1(n576), .A2(n575), .B1(n760), .B2(n574), .ZN(n577) );
  AOI21_X1 U749 ( .B1(n62), .B2(n578), .A(n577), .ZN(n616) );
  OAI22_X1 U750 ( .A1(n579), .A2(n651), .B1(n616), .B2(n797), .ZN(n580) );
  AOI211_X1 U751 ( .C1(n823), .C2(n582), .A(n581), .B(n580), .ZN(n584) );
  OAI211_X1 U752 ( .C1(n585), .C2(n637), .A(n584), .B(n583), .ZN(n598) );
  AOI22_X1 U753 ( .A1(n802), .A2(n587), .B1(n740), .B2(n586), .ZN(n595) );
  AOI22_X1 U754 ( .A1(n62), .A2(n589), .B1(data_in[30]), .B2(n588), .ZN(n590)
         );
  OAI21_X1 U755 ( .B1(n591), .B2(n760), .A(n590), .ZN(n641) );
  AOI22_X1 U756 ( .A1(n810), .A2(n641), .B1(n593), .B2(n592), .ZN(n594) );
  OAI211_X1 U757 ( .C1(n596), .C2(n719), .A(n595), .B(n594), .ZN(n597) );
  AOI211_X1 U758 ( .C1(n634), .C2(n631), .A(n598), .B(n597), .ZN(n599) );
  NAND4_X1 U759 ( .A1(n602), .A2(n601), .A3(n600), .A4(n599), .ZN(data_out[30]) );
  AOI21_X1 U760 ( .B1(n810), .B2(n787), .A(n782), .ZN(n603) );
  AOI221_X1 U761 ( .B1(n606), .B2(n605), .C1(n604), .C2(n605), .A(n603), .ZN(
        n612) );
  AOI21_X1 U762 ( .B1(n807), .B2(n787), .A(n776), .ZN(n609) );
  AOI21_X1 U763 ( .B1(data_in[23]), .B2(n607), .A(n64), .ZN(n608) );
  OAI22_X1 U764 ( .A1(n610), .A2(n834), .B1(n609), .B2(n608), .ZN(n611) );
  OAI22_X1 U765 ( .A1(n616), .A2(n827), .B1(n615), .B2(n614), .ZN(n617) );
  AOI21_X1 U766 ( .B1(n619), .B2(n618), .A(n617), .ZN(n643) );
  AOI22_X1 U767 ( .A1(n623), .A2(n622), .B1(n621), .B2(n620), .ZN(n626) );
  OAI22_X1 U768 ( .A1(n626), .A2(n70), .B1(n625), .B2(n624), .ZN(n640) );
  OAI22_X1 U769 ( .A1(n668), .A2(n629), .B1(n628), .B2(n627), .ZN(n630) );
  INV_X1 U770 ( .A(n630), .ZN(n636) );
  AOI22_X1 U771 ( .A1(n634), .A2(n633), .B1(n632), .B2(n631), .ZN(n635) );
  OAI211_X1 U772 ( .C1(n638), .C2(n637), .A(n636), .B(n635), .ZN(n639) );
  AOI211_X1 U773 ( .C1(n778), .C2(n641), .A(n640), .B(n639), .ZN(n642) );
  OAI22_X1 U774 ( .A1(n646), .A2(n758), .B1(n645), .B2(n757), .ZN(n647) );
  AOI21_X1 U775 ( .B1(n789), .B2(n702), .A(n647), .ZN(n648) );
  OAI21_X1 U776 ( .B1(n705), .B2(n795), .A(n648), .ZN(n685) );
  AOI21_X1 U777 ( .B1(data_in[14]), .B2(n681), .A(n649), .ZN(n698) );
  OAI22_X1 U778 ( .A1(n674), .A2(n651), .B1(n698), .B2(n650), .ZN(n655) );
  OAI22_X1 U779 ( .A1(n653), .A2(n652), .B1(n696), .B2(n678), .ZN(n654) );
  AOI211_X1 U780 ( .C1(n802), .C2(n656), .A(n655), .B(n654), .ZN(n667) );
  INV_X1 U781 ( .A(n657), .ZN(n717) );
  AOI21_X1 U782 ( .B1(n670), .B2(n717), .A(n669), .ZN(n665) );
  AOI21_X1 U783 ( .B1(n716), .B2(n691), .A(n671), .ZN(n664) );
  AOI22_X1 U784 ( .A1(n68), .A2(n761), .B1(n681), .B2(data_in[6]), .ZN(n712)
         );
  OAI22_X1 U785 ( .A1(n712), .A2(n677), .B1(n683), .B2(n743), .ZN(n663) );
  INV_X1 U786 ( .A(n658), .ZN(n659) );
  OAI22_X1 U787 ( .A1(n661), .A2(n660), .B1(n659), .B2(n767), .ZN(n662) );
  NOR4_X1 U788 ( .A1(n665), .A2(n664), .A3(n663), .A4(n662), .ZN(n666) );
  OAI211_X1 U789 ( .C1(n668), .C2(n685), .A(n667), .B(n666), .ZN(data_out[3])
         );
  OAI22_X1 U790 ( .A1(n670), .A2(n715), .B1(n716), .B2(n669), .ZN(n695) );
  OAI22_X1 U791 ( .A1(n712), .A2(n719), .B1(n671), .B2(n717), .ZN(n694) );
  NOR2_X1 U792 ( .A1(n673), .A2(n672), .ZN(n739) );
  INV_X1 U793 ( .A(n674), .ZN(n675) );
  NOR2_X1 U794 ( .A1(n676), .A2(n675), .ZN(n736) );
  OAI22_X1 U795 ( .A1(n739), .A2(n678), .B1(n736), .B2(n677), .ZN(n693) );
  AOI22_X1 U796 ( .A1(n62), .A2(n734), .B1(n679), .B2(n72), .ZN(n722) );
  AOI21_X1 U797 ( .B1(data_in[15]), .B2(n681), .A(n680), .ZN(n728) );
  INV_X1 U798 ( .A(n728), .ZN(n700) );
  AOI22_X1 U799 ( .A1(n823), .A2(n722), .B1(n682), .B2(n700), .ZN(n690) );
  INV_X1 U800 ( .A(n683), .ZN(n688) );
  OAI22_X1 U801 ( .A1(n698), .A2(n684), .B1(n696), .B2(n709), .ZN(n687) );
  OAI22_X1 U802 ( .A1(n834), .A2(n685), .B1(n708), .B2(n743), .ZN(n686) );
  AOI211_X1 U803 ( .C1(n688), .C2(n740), .A(n687), .B(n686), .ZN(n689) );
  OAI211_X1 U804 ( .C1(n718), .C2(n691), .A(n690), .B(n689), .ZN(n692) );
  AOI222_X1 U805 ( .A1(n696), .A2(n62), .B1(n713), .B2(n789), .C1(n787), .C2(
        n711), .ZN(n730) );
  AOI222_X1 U806 ( .A1(n699), .A2(n786), .B1(n72), .B2(n698), .C1(n697), .C2(
        n792), .ZN(n735) );
  AOI22_X1 U807 ( .A1(n810), .A2(n730), .B1(n776), .B2(n735), .ZN(n726) );
  AOI22_X1 U808 ( .A1(n741), .A2(n765), .B1(n701), .B2(n700), .ZN(n725) );
  AOI22_X1 U809 ( .A1(n786), .A2(n703), .B1(n792), .B2(n702), .ZN(n704) );
  OAI21_X1 U810 ( .B1(n705), .B2(n758), .A(n704), .ZN(n706) );
  AOI21_X1 U811 ( .B1(n789), .B2(n707), .A(n706), .ZN(n746) );
  OAI22_X1 U812 ( .A1(n739), .A2(n709), .B1(n708), .B2(n767), .ZN(n710) );
  AOI21_X1 U813 ( .B1(n823), .B2(n746), .A(n710), .ZN(n724) );
  AOI222_X1 U814 ( .A1(n713), .A2(n792), .B1(n712), .B2(n72), .C1(n786), .C2(
        n711), .ZN(n714) );
  INV_X1 U815 ( .A(n714), .ZN(n738) );
  OAI22_X1 U816 ( .A1(n716), .A2(n715), .B1(n818), .B2(n738), .ZN(n721) );
  OAI22_X1 U817 ( .A1(n736), .A2(n719), .B1(n718), .B2(n717), .ZN(n720) );
  AOI211_X1 U818 ( .C1(n802), .C2(n722), .A(n721), .B(n720), .ZN(n723) );
  NAND4_X1 U819 ( .A1(n726), .A2(n725), .A3(n724), .A4(n723), .ZN(data_out[5])
         );
  AOI222_X1 U820 ( .A1(n729), .A2(n792), .B1(n72), .B2(n728), .C1(n727), .C2(
        n786), .ZN(n753) );
  AOI22_X1 U821 ( .A1(n778), .A2(n730), .B1(n776), .B2(n753), .ZN(n749) );
  OAI21_X1 U822 ( .B1(n732), .B2(n731), .A(n62), .ZN(n733) );
  OAI21_X1 U823 ( .B1(n62), .B2(n734), .A(n733), .ZN(n750) );
  AOI22_X1 U824 ( .A1(n823), .A2(n750), .B1(n821), .B2(n735), .ZN(n748) );
  AOI222_X1 U825 ( .A1(n785), .A2(n792), .B1(n736), .B2(n72), .C1(n786), .C2(
        n791), .ZN(n754) );
  INV_X1 U826 ( .A(n754), .ZN(n737) );
  OAI22_X1 U827 ( .A1(n812), .A2(n738), .B1(n818), .B2(n737), .ZN(n745) );
  AOI222_X1 U828 ( .A1(n62), .A2(n739), .B1(n787), .B2(n791), .C1(n789), .C2(
        n785), .ZN(n755) );
  AOI22_X1 U829 ( .A1(n741), .A2(n740), .B1(n810), .B2(n755), .ZN(n742) );
  OAI21_X1 U830 ( .B1(n768), .B2(n743), .A(n742), .ZN(n744) );
  AOI211_X1 U831 ( .C1(n802), .C2(n746), .A(n745), .B(n744), .ZN(n747) );
  NAND3_X1 U832 ( .A1(n749), .A2(n748), .A3(n747), .ZN(data_out[6]) );
  AOI22_X1 U833 ( .A1(n802), .A2(n750), .B1(n776), .B2(n774), .ZN(n773) );
  OAI22_X1 U834 ( .A1(n759), .A2(n757), .B1(n758), .B2(n756), .ZN(n752) );
  OAI22_X1 U835 ( .A1(n795), .A2(n761), .B1(n762), .B2(n760), .ZN(n751) );
  NOR2_X1 U836 ( .A1(n752), .A2(n751), .ZN(n783) );
  AOI22_X1 U837 ( .A1(n782), .A2(n783), .B1(n821), .B2(n753), .ZN(n772) );
  AOI22_X1 U838 ( .A1(n778), .A2(n755), .B1(n784), .B2(n754), .ZN(n771) );
  OAI22_X1 U839 ( .A1(n759), .A2(n758), .B1(n757), .B2(n756), .ZN(n764) );
  OAI22_X1 U840 ( .A1(n795), .A2(n762), .B1(n761), .B2(n760), .ZN(n763) );
  NOR2_X1 U841 ( .A1(n764), .A2(n763), .ZN(n777) );
  AOI22_X1 U842 ( .A1(n64), .A2(n765), .B1(n810), .B2(n777), .ZN(n766) );
  OAI21_X1 U843 ( .B1(n768), .B2(n767), .A(n766), .ZN(n769) );
  AOI21_X1 U844 ( .B1(n823), .B2(n801), .A(n769), .ZN(n770) );
  NAND4_X1 U845 ( .A1(n773), .A2(n772), .A3(n771), .A4(n770), .ZN(data_out[7])
         );
  AOI22_X1 U846 ( .A1(n823), .A2(n775), .B1(n821), .B2(n774), .ZN(n806) );
  AOI22_X1 U847 ( .A1(n778), .A2(n777), .B1(n820), .B2(n776), .ZN(n805) );
  AOI22_X1 U848 ( .A1(n788), .A2(n786), .B1(n787), .B2(n785), .ZN(n780) );
  AOI22_X1 U849 ( .A1(n792), .A2(n790), .B1(n791), .B2(n789), .ZN(n779) );
  NAND2_X1 U850 ( .A1(n780), .A2(n779), .ZN(n811) );
  INV_X1 U851 ( .A(n811), .ZN(n781) );
  AOI22_X1 U852 ( .A1(n784), .A2(n783), .B1(n782), .B2(n781), .ZN(n804) );
  AOI22_X1 U853 ( .A1(n788), .A2(n787), .B1(n786), .B2(n785), .ZN(n794) );
  AOI22_X1 U854 ( .A1(n792), .A2(n791), .B1(n790), .B2(n789), .ZN(n793) );
  NAND2_X1 U855 ( .A1(n794), .A2(n793), .ZN(n813) );
  NAND2_X1 U856 ( .A1(n796), .A2(n795), .ZN(n826) );
  OAI22_X1 U857 ( .A1(n798), .A2(n813), .B1(n797), .B2(n826), .ZN(n799) );
  AOI211_X1 U858 ( .C1(n802), .C2(n801), .A(n800), .B(n799), .ZN(n803) );
  NAND4_X1 U859 ( .A1(n806), .A2(n805), .A3(n804), .A4(n803), .ZN(data_out[8])
         );
  AOI22_X1 U860 ( .A1(n810), .A2(n809), .B1(n808), .B2(n807), .ZN(n832) );
  OAI22_X1 U861 ( .A1(n814), .A2(n813), .B1(n812), .B2(n811), .ZN(n830) );
  INV_X1 U862 ( .A(n815), .ZN(n817) );
  OAI22_X1 U863 ( .A1(n819), .A2(n818), .B1(n817), .B2(n816), .ZN(n829) );
  AOI22_X1 U864 ( .A1(n823), .A2(n822), .B1(n821), .B2(n820), .ZN(n825) );
  OAI211_X1 U865 ( .C1(n827), .C2(n826), .A(n825), .B(n824), .ZN(n828) );
  NOR3_X1 U866 ( .A1(n830), .A2(n829), .A3(n828), .ZN(n831) );
  OAI211_X1 U867 ( .C1(n834), .C2(n833), .A(n832), .B(n831), .ZN(data_out[9])
         );
endmodule


module a_generator ( a_in, neg_a_in, sel, a, neg_a, ax2, neg_ax2 );
  input [63:0] a_in;
  input [63:0] neg_a_in;
  input [3:0] sel;
  output [63:0] a;
  output [63:0] neg_a;
  output [63:0] ax2;
  output [63:0] neg_ax2;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736;

  INV_X1 U2 ( .A(n574), .ZN(n1) );
  NAND2_X1 U3 ( .A1(n539), .A2(n589), .ZN(n2) );
  OAI21_X1 U4 ( .B1(n103), .B2(n547), .A(n2), .ZN(n3) );
  OAI22_X1 U5 ( .A1(n93), .A2(n517), .B1(n100), .B2(n516), .ZN(n4) );
  AOI211_X1 U6 ( .C1(n126), .C2(n518), .A(n3), .B(n4), .ZN(n5) );
  OAI21_X1 U7 ( .B1(n91), .B2(n1), .A(n5), .ZN(a[30]) );
  AOI22_X1 U8 ( .A1(n723), .A2(a_in[53]), .B1(n128), .B2(a_in[27]), .ZN(n6) );
  AOI22_X1 U9 ( .A1(n114), .A2(a_in[49]), .B1(n130), .B2(a_in[55]), .ZN(n7) );
  AOI22_X1 U10 ( .A1(n92), .A2(a_in[51]), .B1(n122), .B2(n698), .ZN(n8) );
  AOI22_X1 U11 ( .A1(n700), .A2(n717), .B1(n118), .B2(n699), .ZN(n9) );
  AND4_X1 U12 ( .A1(n6), .A2(n7), .A3(n8), .A4(n9), .ZN(n10) );
  OAI21_X1 U13 ( .B1(n97), .B2(n679), .A(n10), .ZN(a[57]) );
  INV_X1 U14 ( .A(n278), .ZN(n11) );
  NAND2_X1 U15 ( .A1(n539), .A2(n295), .ZN(n12) );
  OAI21_X1 U16 ( .B1(n103), .B2(n248), .A(n12), .ZN(n13) );
  OAI22_X1 U17 ( .A1(n93), .A2(n229), .B1(n100), .B2(n228), .ZN(n14) );
  AOI211_X1 U18 ( .C1(n126), .C2(n230), .A(n13), .B(n14), .ZN(n15) );
  OAI21_X1 U19 ( .B1(n119), .B2(n11), .A(n15), .ZN(neg_a[31]) );
  AOI22_X1 U20 ( .A1(n723), .A2(neg_a_in[55]), .B1(n128), .B2(neg_a_in[29]), 
        .ZN(n16) );
  AOI22_X1 U21 ( .A1(n114), .A2(neg_a_in[51]), .B1(n129), .B2(neg_a_in[57]), 
        .ZN(n17) );
  AOI22_X1 U22 ( .A1(n92), .A2(neg_a_in[53]), .B1(n122), .B2(n712), .ZN(n18)
         );
  AOI22_X1 U23 ( .A1(n713), .A2(n717), .B1(n118), .B2(n714), .ZN(n19) );
  AND4_X1 U24 ( .A1(n16), .A2(n17), .A3(n18), .A4(n19), .ZN(n20) );
  OAI21_X1 U25 ( .B1(n97), .B2(n386), .A(n20), .ZN(neg_a[59]) );
  AOI22_X1 U26 ( .A1(n114), .A2(neg_a_in[4]), .B1(neg_a_in[8]), .B2(n723), 
        .ZN(n21) );
  AOI22_X1 U27 ( .A1(n129), .A2(neg_a_in[10]), .B1(neg_a_in[6]), .B2(n92), 
        .ZN(n22) );
  AOI22_X1 U28 ( .A1(n724), .A2(neg_a_in[0]), .B1(n95), .B2(neg_a_in[2]), .ZN(
        n23) );
  NAND3_X1 U29 ( .A1(n21), .A2(n22), .A3(n23), .ZN(neg_a[12]) );
  INV_X1 U30 ( .A(n282), .ZN(n24) );
  NAND2_X1 U31 ( .A1(n539), .A2(n283), .ZN(n25) );
  OAI21_X1 U32 ( .B1(n103), .B2(n257), .A(n25), .ZN(n26) );
  OAI22_X1 U33 ( .A1(n93), .A2(n233), .B1(n100), .B2(n232), .ZN(n27) );
  AOI211_X1 U34 ( .C1(n126), .C2(n234), .A(n26), .B(n27), .ZN(n28) );
  OAI21_X1 U35 ( .B1(n119), .B2(n24), .A(n28), .ZN(neg_a[32]) );
  AOI22_X1 U36 ( .A1(n723), .A2(a_in[52]), .B1(n128), .B2(a_in[26]), .ZN(n29)
         );
  AOI22_X1 U37 ( .A1(n114), .A2(a_in[48]), .B1(n129), .B2(a_in[54]), .ZN(n30)
         );
  AOI22_X1 U38 ( .A1(n92), .A2(a_in[50]), .B1(n122), .B2(n688), .ZN(n31) );
  AOI22_X1 U39 ( .A1(n690), .A2(n717), .B1(n118), .B2(n689), .ZN(n32) );
  AND4_X1 U40 ( .A1(n29), .A2(n30), .A3(n31), .A4(n32), .ZN(n33) );
  OAI21_X1 U41 ( .B1(n97), .B2(n678), .A(n33), .ZN(a[56]) );
  INV_X1 U42 ( .A(n287), .ZN(n34) );
  NAND2_X1 U43 ( .A1(n539), .A2(n288), .ZN(n35) );
  OAI21_X1 U44 ( .B1(n103), .B2(n266), .A(n35), .ZN(n36) );
  OAI22_X1 U45 ( .A1(n93), .A2(n237), .B1(n100), .B2(n236), .ZN(n37) );
  AOI211_X1 U46 ( .C1(n126), .C2(n238), .A(n36), .B(n37), .ZN(n38) );
  OAI21_X1 U47 ( .B1(n119), .B2(n34), .A(n38), .ZN(neg_a[33]) );
  NAND3_X1 U48 ( .A1(n109), .A2(n133), .A3(neg_a_in[4]), .ZN(n39) );
  NAND2_X1 U49 ( .A1(n497), .A2(neg_a_in[2]), .ZN(n40) );
  OAI211_X1 U50 ( .C1(n109), .C2(n242), .A(n39), .B(n40), .ZN(n223) );
  AOI22_X1 U51 ( .A1(n723), .A2(neg_a_in[54]), .B1(neg_a_in[28]), .B2(n128), 
        .ZN(n41) );
  AOI22_X1 U52 ( .A1(n114), .A2(neg_a_in[50]), .B1(n130), .B2(neg_a_in[56]), 
        .ZN(n42) );
  AOI22_X1 U53 ( .A1(n92), .A2(neg_a_in[52]), .B1(n122), .B2(n410), .ZN(n43)
         );
  AOI22_X1 U54 ( .A1(n411), .A2(n717), .B1(n118), .B2(n412), .ZN(n44) );
  AND4_X1 U55 ( .A1(n41), .A2(n42), .A3(n43), .A4(n44), .ZN(n45) );
  OAI21_X1 U56 ( .B1(n97), .B2(n385), .A(n45), .ZN(neg_a[58]) );
  INV_X1 U57 ( .A(n103), .ZN(n46) );
  INV_X1 U58 ( .A(n100), .ZN(n47) );
  AOI222_X1 U59 ( .A1(n46), .A2(n407), .B1(n94), .B2(n378), .C1(n47), .C2(
        neg_a_in[23]), .ZN(n48) );
  OR2_X1 U60 ( .A1(n358), .A2(n124), .ZN(n49) );
  OAI211_X1 U61 ( .C1(n93), .C2(n379), .A(n48), .B(n49), .ZN(neg_a[53]) );
  AOI22_X1 U62 ( .A1(n723), .A2(a_in[55]), .B1(n128), .B2(a_in[29]), .ZN(n50)
         );
  AOI22_X1 U63 ( .A1(n114), .A2(a_in[51]), .B1(n130), .B2(a_in[57]), .ZN(n51)
         );
  AOI22_X1 U64 ( .A1(n92), .A2(a_in[53]), .B1(n122), .B2(n715), .ZN(n52) );
  AOI22_X1 U65 ( .A1(n720), .A2(n717), .B1(n118), .B2(n716), .ZN(n53) );
  AND4_X1 U66 ( .A1(n50), .A2(n51), .A3(n52), .A4(n53), .ZN(n54) );
  OAI21_X1 U67 ( .B1(n97), .B2(n687), .A(n54), .ZN(a[59]) );
  AOI22_X1 U68 ( .A1(n497), .A2(neg_a_in[5]), .B1(n498), .B2(neg_a_in[7]), 
        .ZN(n55) );
  OAI21_X1 U69 ( .B1(n109), .B2(n268), .A(n55), .ZN(n238) );
  AOI22_X1 U70 ( .A1(n721), .A2(n411), .B1(n118), .B2(n410), .ZN(n56) );
  AOI22_X1 U71 ( .A1(n129), .A2(neg_a_in[60]), .B1(n128), .B2(neg_a_in[32]), 
        .ZN(n57) );
  AOI22_X1 U72 ( .A1(n95), .A2(neg_a_in[52]), .B1(n412), .B2(n717), .ZN(n58)
         );
  AOI22_X1 U73 ( .A1(n92), .A2(neg_a_in[56]), .B1(n723), .B2(neg_a_in[58]), 
        .ZN(n59) );
  AND4_X1 U74 ( .A1(n56), .A2(n57), .A3(n58), .A4(n59), .ZN(n60) );
  AOI22_X1 U75 ( .A1(n724), .A2(neg_a_in[50]), .B1(n114), .B2(neg_a_in[54]), 
        .ZN(n61) );
  AOI22_X1 U76 ( .A1(n726), .A2(neg_a_in[46]), .B1(n725), .B2(neg_a_in[48]), 
        .ZN(n62) );
  NAND3_X1 U77 ( .A1(n60), .A2(n61), .A3(n62), .ZN(neg_a[62]) );
  AOI22_X1 U78 ( .A1(n497), .A2(neg_a_in[4]), .B1(n498), .B2(neg_a_in[6]), 
        .ZN(n63) );
  OAI21_X1 U79 ( .B1(n109), .B2(n259), .A(n63), .ZN(n234) );
  AOI22_X1 U80 ( .A1(n717), .A2(n710), .B1(n118), .B2(n709), .ZN(n64) );
  AOI22_X1 U81 ( .A1(n130), .A2(a_in[60]), .B1(n128), .B2(a_in[32]), .ZN(n65)
         );
  AOI22_X1 U82 ( .A1(n95), .A2(a_in[52]), .B1(n711), .B2(n721), .ZN(n66) );
  AOI22_X1 U83 ( .A1(n92), .A2(a_in[56]), .B1(n723), .B2(a_in[58]), .ZN(n67)
         );
  AND4_X1 U84 ( .A1(n64), .A2(n65), .A3(n66), .A4(n67), .ZN(n68) );
  AOI22_X1 U85 ( .A1(n724), .A2(a_in[50]), .B1(n114), .B2(a_in[54]), .ZN(n69)
         );
  AOI22_X1 U86 ( .A1(n725), .A2(a_in[48]), .B1(n726), .B2(a_in[46]), .ZN(n70)
         );
  NAND3_X1 U87 ( .A1(n68), .A2(n69), .A3(n70), .ZN(a[62]) );
  AOI22_X1 U88 ( .A1(n717), .A2(n716), .B1(n118), .B2(n715), .ZN(n71) );
  AOI22_X1 U89 ( .A1(n130), .A2(a_in[61]), .B1(n128), .B2(a_in[33]), .ZN(n72)
         );
  AOI22_X1 U90 ( .A1(n95), .A2(a_in[53]), .B1(n720), .B2(n721), .ZN(n73) );
  AOI22_X1 U91 ( .A1(n92), .A2(a_in[57]), .B1(n723), .B2(a_in[59]), .ZN(n74)
         );
  AND4_X1 U92 ( .A1(n71), .A2(n72), .A3(n73), .A4(n74), .ZN(n75) );
  AOI22_X1 U93 ( .A1(n724), .A2(a_in[51]), .B1(n114), .B2(a_in[55]), .ZN(n76)
         );
  AOI22_X1 U94 ( .A1(n725), .A2(a_in[49]), .B1(n726), .B2(a_in[47]), .ZN(n77)
         );
  NAND3_X1 U95 ( .A1(n75), .A2(n76), .A3(n77), .ZN(a[63]) );
  AOI22_X1 U96 ( .A1(n713), .A2(n721), .B1(n118), .B2(n712), .ZN(n78) );
  AOI22_X1 U97 ( .A1(n130), .A2(neg_a_in[61]), .B1(n128), .B2(neg_a_in[33]), 
        .ZN(n79) );
  AOI22_X1 U98 ( .A1(n95), .A2(neg_a_in[53]), .B1(n717), .B2(n714), .ZN(n80)
         );
  AOI22_X1 U99 ( .A1(n92), .A2(neg_a_in[57]), .B1(n723), .B2(neg_a_in[59]), 
        .ZN(n81) );
  AND4_X1 U100 ( .A1(n78), .A2(n79), .A3(n80), .A4(n81), .ZN(n82) );
  AOI22_X1 U101 ( .A1(n724), .A2(neg_a_in[51]), .B1(n114), .B2(neg_a_in[55]), 
        .ZN(n83) );
  AOI22_X1 U102 ( .A1(n725), .A2(neg_a_in[49]), .B1(n726), .B2(neg_a_in[47]), 
        .ZN(n84) );
  NAND3_X1 U103 ( .A1(n82), .A2(n83), .A3(n84), .ZN(neg_a[63]) );
  AND2_X4 U104 ( .A1(n98), .A2(n113), .ZN(n114) );
  INV_X2 U105 ( .A(n722), .ZN(n92) );
  INV_X4 U106 ( .A(n116), .ZN(n723) );
  INV_X2 U107 ( .A(n718), .ZN(n130) );
  INV_X2 U108 ( .A(n718), .ZN(n129) );
  BUF_X1 U109 ( .A(n136), .Z(n85) );
  BUF_X2 U110 ( .A(n136), .Z(n86) );
  INV_X1 U111 ( .A(sel[3]), .ZN(n136) );
  OR2_X2 U112 ( .A1(n644), .A2(n120), .ZN(n116) );
  OR2_X2 U113 ( .A1(n87), .A2(n120), .ZN(n115) );
  CLKBUF_X3 U114 ( .A(n644), .Z(n87) );
  AND2_X2 U115 ( .A1(n127), .A2(n98), .ZN(n724) );
  INV_X2 U116 ( .A(n724), .ZN(n465) );
  CLKBUF_X3 U117 ( .A(n643), .Z(n88) );
  NAND2_X1 U118 ( .A1(n86), .A2(n106), .ZN(n103) );
  OR2_X1 U119 ( .A1(n218), .A2(n135), .ZN(n100) );
  INV_X1 U120 ( .A(n133), .ZN(n89) );
  INV_X1 U121 ( .A(n87), .ZN(n98) );
  INV_X1 U122 ( .A(n93), .ZN(n90) );
  INV_X1 U123 ( .A(n94), .ZN(n91) );
  INV_X1 U124 ( .A(sel[0]), .ZN(n133) );
  BUF_X1 U125 ( .A(n719), .Z(n95) );
  INV_X1 U126 ( .A(n126), .ZN(n97) );
  NAND2_X1 U127 ( .A1(n85), .A2(sel[0]), .ZN(n644) );
  INV_X2 U128 ( .A(n113), .ZN(n93) );
  INV_X2 U129 ( .A(n133), .ZN(n132) );
  BUF_X2 U130 ( .A(n605), .Z(n94) );
  OR2_X1 U131 ( .A1(sel[3]), .A2(sel[0]), .ZN(n643) );
  INV_X1 U132 ( .A(n114), .ZN(n96) );
  INV_X1 U133 ( .A(n126), .ZN(n124) );
  NAND2_X2 U134 ( .A1(n329), .A2(n605), .ZN(n718) );
  NAND2_X1 U135 ( .A1(n329), .A2(n113), .ZN(n722) );
  BUF_X1 U136 ( .A(n86), .Z(n135) );
  INV_X1 U137 ( .A(n133), .ZN(n111) );
  INV_X4 U138 ( .A(n103), .ZN(n122) );
  INV_X4 U139 ( .A(n100), .ZN(n128) );
  INV_X2 U140 ( .A(n86), .ZN(n134) );
  AND2_X1 U141 ( .A1(n90), .A2(n135), .ZN(n539) );
  INV_X1 U142 ( .A(n719), .ZN(n464) );
  AND2_X1 U143 ( .A1(n123), .A2(n132), .ZN(n726) );
  NOR2_X1 U144 ( .A1(n125), .A2(n88), .ZN(n719) );
  INV_X1 U145 ( .A(n507), .ZN(n497) );
  NAND2_X1 U146 ( .A1(n109), .A2(n131), .ZN(n507) );
  INV_X1 U147 ( .A(n133), .ZN(n131) );
  INV_X1 U148 ( .A(n440), .ZN(n486) );
  INV_X1 U149 ( .A(n127), .ZN(n125) );
  NOR2_X1 U150 ( .A1(n110), .A2(sel[1]), .ZN(n127) );
  INV_X1 U151 ( .A(sel[2]), .ZN(n110) );
  INV_X1 U152 ( .A(sel[1]), .ZN(n141) );
  INV_X1 U153 ( .A(n510), .ZN(n498) );
  OR2_X1 U154 ( .A1(n86), .A2(n89), .ZN(n510) );
  INV_X1 U155 ( .A(n134), .ZN(n112) );
  AND2_X1 U156 ( .A1(n123), .A2(n133), .ZN(n725) );
  INV_X1 U157 ( .A(n439), .ZN(n485) );
  AND2_X1 U158 ( .A1(n121), .A2(n134), .ZN(n717) );
  AND2_X1 U159 ( .A1(n94), .A2(n134), .ZN(n118) );
  INV_X1 U160 ( .A(n86), .ZN(n109) );
  BUF_X2 U161 ( .A(n127), .Z(n126) );
  INV_X2 U162 ( .A(n93), .ZN(n121) );
  INV_X2 U163 ( .A(n94), .ZN(n119) );
  OAI21_X1 U164 ( .B1(n397), .B2(n125), .A(n396), .ZN(neg_a[60]) );
  AOI211_X1 U165 ( .C1(n395), .C2(n717), .A(n394), .B(n393), .ZN(n396) );
  OAI21_X1 U166 ( .B1(n96), .B2(n392), .A(n391), .ZN(n393) );
  AOI22_X1 U167 ( .A1(n723), .A2(neg_a_in[56]), .B1(neg_a_in[30]), .B2(n128), 
        .ZN(n391) );
  OAI211_X1 U168 ( .C1(n402), .C2(n390), .A(n389), .B(n388), .ZN(n394) );
  AOI22_X1 U169 ( .A1(n92), .A2(neg_a_in[54]), .B1(n130), .B2(neg_a_in[58]), 
        .ZN(n388) );
  INV_X1 U170 ( .A(neg_a_in[44]), .ZN(n390) );
  NAND4_X1 U171 ( .A1(n99), .A2(n697), .A3(n696), .A4(n695), .ZN(a[60]) );
  AOI22_X1 U172 ( .A1(n723), .A2(a_in[56]), .B1(n92), .B2(a_in[54]), .ZN(n697)
         );
  NAND2_X1 U173 ( .A1(n721), .A2(n690), .ZN(n691) );
  NAND2_X1 U174 ( .A1(n95), .A2(a_in[50]), .ZN(n692) );
  AOI22_X1 U175 ( .A1(n130), .A2(a_in[58]), .B1(n128), .B2(a_in[30]), .ZN(n693) );
  AOI22_X1 U176 ( .A1(n717), .A2(n689), .B1(n118), .B2(n688), .ZN(n694) );
  OAI211_X1 U177 ( .C1(n686), .C2(n125), .A(n685), .B(n684), .ZN(a[58]) );
  AOI22_X1 U178 ( .A1(n717), .A2(n711), .B1(n118), .B2(n710), .ZN(n684) );
  AND4_X1 U179 ( .A1(n683), .A2(n682), .A3(n681), .A4(n680), .ZN(n685) );
  NAND2_X1 U180 ( .A1(n709), .A2(n122), .ZN(n680) );
  NAND2_X1 U181 ( .A1(n92), .A2(a_in[52]), .ZN(n681) );
  AOI22_X1 U182 ( .A1(n723), .A2(a_in[54]), .B1(n128), .B2(a_in[28]), .ZN(n682) );
  NAND4_X1 U183 ( .A1(n708), .A2(n707), .A3(n706), .A4(n705), .ZN(a[61]) );
  AOI22_X1 U184 ( .A1(n723), .A2(a_in[57]), .B1(n92), .B2(a_in[55]), .ZN(n707)
         );
  AND4_X1 U185 ( .A1(n704), .A2(n703), .A3(n702), .A4(n701), .ZN(n708) );
  NAND2_X1 U186 ( .A1(n721), .A2(n700), .ZN(n701) );
  NAND2_X1 U187 ( .A1(n95), .A2(a_in[51]), .ZN(n702) );
  AOI22_X1 U188 ( .A1(n130), .A2(a_in[59]), .B1(n128), .B2(a_in[31]), .ZN(n703) );
  AOI22_X1 U189 ( .A1(n717), .A2(n699), .B1(n118), .B2(n698), .ZN(n704) );
  OAI21_X1 U190 ( .B1(n409), .B2(n125), .A(n408), .ZN(neg_a[61]) );
  AOI211_X1 U191 ( .C1(n407), .C2(n717), .A(n406), .B(n405), .ZN(n408) );
  OAI21_X1 U192 ( .B1(n96), .B2(n404), .A(n403), .ZN(n405) );
  AOI22_X1 U193 ( .A1(n723), .A2(neg_a_in[57]), .B1(n128), .B2(neg_a_in[31]), 
        .ZN(n403) );
  OAI211_X1 U194 ( .C1(n402), .C2(n401), .A(n400), .B(n399), .ZN(n406) );
  INV_X1 U195 ( .A(neg_a_in[45]), .ZN(n401) );
  INV_X1 U196 ( .A(n726), .ZN(n402) );
  NOR2_X1 U197 ( .A1(n125), .A2(n112), .ZN(n721) );
  OAI21_X1 U198 ( .B1(n409), .B2(n93), .A(n384), .ZN(neg_a[57]) );
  AOI21_X1 U199 ( .B1(n383), .B2(n126), .A(n382), .ZN(n384) );
  AOI22_X1 U200 ( .A1(n129), .A2(neg_a_in[55]), .B1(n128), .B2(neg_a_in[27]), 
        .ZN(n380) );
  AOI22_X1 U201 ( .A1(n118), .A2(n407), .B1(n398), .B2(n122), .ZN(n381) );
  INV_X1 U202 ( .A(neg_a_in[53]), .ZN(n404) );
  INV_X1 U203 ( .A(n379), .ZN(n383) );
  OAI21_X1 U204 ( .B1(n677), .B2(n124), .A(n676), .ZN(a[55]) );
  AOI21_X1 U205 ( .B1(n675), .B2(n90), .A(n674), .ZN(n676) );
  AOI22_X1 U206 ( .A1(n130), .A2(a_in[53]), .B1(n128), .B2(a_in[25]), .ZN(n671) );
  AOI22_X1 U207 ( .A1(n118), .A2(n720), .B1(n716), .B2(n122), .ZN(n672) );
  INV_X1 U208 ( .A(a_in[51]), .ZN(n673) );
  INV_X1 U209 ( .A(n687), .ZN(n675) );
  OAI21_X1 U210 ( .B1(n370), .B2(n125), .A(n369), .ZN(neg_a[55]) );
  AOI21_X1 U211 ( .B1(n368), .B2(n121), .A(n367), .ZN(n369) );
  AOI22_X1 U212 ( .A1(n129), .A2(neg_a_in[53]), .B1(n128), .B2(neg_a_in[25]), 
        .ZN(n365) );
  AOI22_X1 U213 ( .A1(n118), .A2(n713), .B1(n714), .B2(n122), .ZN(n366) );
  INV_X1 U214 ( .A(n386), .ZN(n368) );
  OAI21_X1 U215 ( .B1(n397), .B2(n93), .A(n377), .ZN(neg_a[56]) );
  AOI21_X1 U216 ( .B1(n376), .B2(n126), .A(n375), .ZN(n377) );
  AOI22_X1 U217 ( .A1(n130), .A2(neg_a_in[54]), .B1(n128), .B2(neg_a_in[26]), 
        .ZN(n373) );
  AOI22_X1 U218 ( .A1(n118), .A2(n395), .B1(n387), .B2(n122), .ZN(n374) );
  INV_X1 U219 ( .A(neg_a_in[52]), .ZN(n392) );
  INV_X1 U220 ( .A(n372), .ZN(n376) );
  OAI21_X1 U221 ( .B1(n364), .B2(n124), .A(n363), .ZN(neg_a[54]) );
  AOI21_X1 U222 ( .B1(n362), .B2(n121), .A(n361), .ZN(n363) );
  AOI22_X1 U223 ( .A1(n130), .A2(neg_a_in[52]), .B1(n128), .B2(neg_a_in[24]), 
        .ZN(n359) );
  AOI22_X1 U224 ( .A1(n118), .A2(n411), .B1(n412), .B2(n122), .ZN(n360) );
  INV_X1 U225 ( .A(n385), .ZN(n362) );
  OAI21_X1 U226 ( .B1(n670), .B2(n124), .A(n669), .ZN(a[54]) );
  AOI21_X1 U227 ( .B1(n668), .B2(n90), .A(n667), .ZN(n669) );
  AOI22_X1 U228 ( .A1(n130), .A2(a_in[52]), .B1(n128), .B2(a_in[24]), .ZN(n664) );
  AOI22_X1 U229 ( .A1(n118), .A2(n711), .B1(n710), .B2(n122), .ZN(n665) );
  INV_X1 U230 ( .A(a_in[50]), .ZN(n666) );
  INV_X1 U231 ( .A(n686), .ZN(n668) );
  OAI21_X1 U232 ( .B1(n663), .B2(n124), .A(n662), .ZN(a[53]) );
  AOI22_X1 U233 ( .A1(n130), .A2(a_in[51]), .B1(n128), .B2(a_in[23]), .ZN(n658) );
  AOI22_X1 U234 ( .A1(n118), .A2(n700), .B1(n699), .B2(n122), .ZN(n659) );
  OAI21_X1 U235 ( .B1(n657), .B2(n124), .A(n656), .ZN(a[52]) );
  AOI22_X1 U236 ( .A1(n130), .A2(a_in[50]), .B1(n128), .B2(a_in[22]), .ZN(n652) );
  AOI22_X1 U237 ( .A1(n118), .A2(n690), .B1(n689), .B2(n122), .ZN(n653) );
  OAI21_X1 U238 ( .B1(n356), .B2(n125), .A(n355), .ZN(neg_a[52]) );
  NOR2_X1 U239 ( .A1(n372), .A2(n93), .ZN(n353) );
  OAI22_X1 U240 ( .A1(n103), .A2(n352), .B1(n100), .B2(n351), .ZN(n354) );
  INV_X1 U241 ( .A(neg_a_in[22]), .ZN(n351) );
  INV_X1 U242 ( .A(n395), .ZN(n352) );
  OAI21_X1 U243 ( .B1(n651), .B2(n124), .A(n650), .ZN(a[51]) );
  AOI21_X1 U244 ( .B1(n121), .B2(n649), .A(n648), .ZN(n650) );
  OAI21_X1 U245 ( .B1(n687), .B2(n119), .A(n647), .ZN(n648) );
  AOI22_X1 U246 ( .A1(n122), .A2(n720), .B1(n128), .B2(a_in[21]), .ZN(n647) );
  AOI21_X1 U247 ( .B1(n646), .B2(n109), .A(n645), .ZN(n687) );
  INV_X1 U248 ( .A(n642), .ZN(n651) );
  OAI21_X1 U249 ( .B1(n349), .B2(n124), .A(n348), .ZN(neg_a[51]) );
  AOI21_X1 U250 ( .B1(n121), .B2(n347), .A(n346), .ZN(n348) );
  OAI21_X1 U251 ( .B1(n386), .B2(n91), .A(n345), .ZN(n346) );
  AOI22_X1 U252 ( .A1(n122), .A2(n713), .B1(n128), .B2(neg_a_in[21]), .ZN(n345) );
  AOI21_X1 U253 ( .B1(n344), .B2(n109), .A(n343), .ZN(n386) );
  INV_X1 U254 ( .A(n342), .ZN(n349) );
  OAI21_X1 U255 ( .B1(n341), .B2(n124), .A(n340), .ZN(neg_a[50]) );
  AOI21_X1 U256 ( .B1(n121), .B2(n339), .A(n338), .ZN(n340) );
  OAI21_X1 U257 ( .B1(n385), .B2(n119), .A(n337), .ZN(n338) );
  AOI22_X1 U258 ( .A1(n122), .A2(n411), .B1(n128), .B2(neg_a_in[20]), .ZN(n337) );
  AOI21_X1 U259 ( .B1(n336), .B2(n109), .A(n335), .ZN(n385) );
  INV_X1 U260 ( .A(n334), .ZN(n341) );
  OAI21_X1 U261 ( .B1(n641), .B2(n125), .A(n640), .ZN(a[50]) );
  AOI21_X1 U262 ( .B1(n121), .B2(n639), .A(n638), .ZN(n640) );
  OAI21_X1 U263 ( .B1(n686), .B2(n119), .A(n637), .ZN(n638) );
  AOI22_X1 U264 ( .A1(n122), .A2(n711), .B1(n128), .B2(a_in[20]), .ZN(n637) );
  AOI21_X1 U265 ( .B1(n636), .B2(n109), .A(n635), .ZN(n686) );
  INV_X1 U266 ( .A(n634), .ZN(n641) );
  OAI21_X1 U267 ( .B1(n358), .B2(n93), .A(n333), .ZN(neg_a[49]) );
  AOI211_X1 U268 ( .C1(n126), .C2(n332), .A(n331), .B(n330), .ZN(n333) );
  NOR2_X1 U269 ( .A1(n379), .A2(n119), .ZN(n330) );
  OAI22_X1 U270 ( .A1(n100), .A2(n327), .B1(n103), .B2(n357), .ZN(n331) );
  OAI21_X1 U271 ( .B1(n663), .B2(n93), .A(n633), .ZN(a[49]) );
  AOI21_X1 U272 ( .B1(n126), .B2(n632), .A(n631), .ZN(n633) );
  OAI21_X1 U273 ( .B1(n679), .B2(n119), .A(n630), .ZN(n631) );
  AOI22_X1 U274 ( .A1(n122), .A2(n700), .B1(n128), .B2(a_in[19]), .ZN(n630) );
  INV_X1 U275 ( .A(a_in[45]), .ZN(n629) );
  INV_X1 U276 ( .A(n627), .ZN(n663) );
  OAI21_X1 U277 ( .B1(n356), .B2(n93), .A(n326), .ZN(neg_a[48]) );
  AOI211_X1 U278 ( .C1(n126), .C2(n325), .A(n324), .B(n323), .ZN(n326) );
  NOR2_X1 U279 ( .A1(n372), .A2(n119), .ZN(n323) );
  OAI22_X1 U280 ( .A1(n100), .A2(n321), .B1(n103), .B2(n350), .ZN(n324) );
  OAI21_X1 U281 ( .B1(n657), .B2(n93), .A(n626), .ZN(a[48]) );
  AOI21_X1 U282 ( .B1(n126), .B2(n625), .A(n624), .ZN(n626) );
  OAI21_X1 U283 ( .B1(n678), .B2(n91), .A(n623), .ZN(n624) );
  AOI22_X1 U284 ( .A1(n122), .A2(n690), .B1(n128), .B2(a_in[18]), .ZN(n623) );
  INV_X1 U285 ( .A(a_in[44]), .ZN(n622) );
  INV_X1 U286 ( .A(n620), .ZN(n657) );
  OAI211_X1 U287 ( .C1(n677), .C2(n91), .A(n619), .B(n618), .ZN(a[47]) );
  AOI22_X1 U288 ( .A1(n646), .A2(n122), .B1(n128), .B2(a_in[17]), .ZN(n618) );
  INV_X1 U289 ( .A(n617), .ZN(n646) );
  AOI22_X1 U290 ( .A1(n126), .A2(n616), .B1(n642), .B2(n121), .ZN(n619) );
  INV_X1 U291 ( .A(n649), .ZN(n677) );
  OAI211_X1 U292 ( .C1(n370), .C2(n91), .A(n320), .B(n319), .ZN(neg_a[47]) );
  AOI22_X1 U293 ( .A1(n344), .A2(n122), .B1(n128), .B2(neg_a_in[17]), .ZN(n319) );
  INV_X1 U294 ( .A(n318), .ZN(n344) );
  AOI22_X1 U295 ( .A1(n126), .A2(n317), .B1(n342), .B2(n121), .ZN(n320) );
  INV_X1 U296 ( .A(n347), .ZN(n370) );
  OAI211_X1 U297 ( .C1(n670), .C2(n119), .A(n614), .B(n613), .ZN(a[46]) );
  AOI22_X1 U298 ( .A1(n636), .A2(n122), .B1(n128), .B2(a_in[16]), .ZN(n613) );
  INV_X1 U299 ( .A(n612), .ZN(n636) );
  AOI22_X1 U300 ( .A1(n126), .A2(n611), .B1(n634), .B2(n121), .ZN(n614) );
  INV_X1 U301 ( .A(n639), .ZN(n670) );
  OAI211_X1 U302 ( .C1(n364), .C2(n91), .A(n315), .B(n314), .ZN(neg_a[46]) );
  AOI22_X1 U303 ( .A1(n336), .A2(n122), .B1(neg_a_in[16]), .B2(n128), .ZN(n314) );
  INV_X1 U304 ( .A(n313), .ZN(n336) );
  AOI22_X1 U305 ( .A1(n126), .A2(n312), .B1(n334), .B2(n121), .ZN(n315) );
  INV_X1 U306 ( .A(n339), .ZN(n364) );
  OAI211_X1 U307 ( .C1(n310), .C2(n97), .A(n309), .B(n308), .ZN(neg_a[45]) );
  AOI22_X1 U308 ( .A1(n122), .A2(n328), .B1(n128), .B2(neg_a_in[15]), .ZN(n308) );
  INV_X1 U309 ( .A(n358), .ZN(n307) );
  INV_X1 U310 ( .A(n398), .ZN(n306) );
  OAI211_X1 U311 ( .C1(n609), .C2(n97), .A(n608), .B(n607), .ZN(a[45]) );
  AOI22_X1 U312 ( .A1(n606), .A2(n122), .B1(n128), .B2(a_in[15]), .ZN(n607) );
  INV_X1 U313 ( .A(n628), .ZN(n606) );
  AOI22_X1 U314 ( .A1(n94), .A2(n627), .B1(n632), .B2(n121), .ZN(n608) );
  INV_X1 U315 ( .A(n603), .ZN(n609) );
  OAI211_X1 U316 ( .C1(n304), .C2(n97), .A(n303), .B(n302), .ZN(neg_a[44]) );
  AOI22_X1 U317 ( .A1(n122), .A2(n322), .B1(n128), .B2(neg_a_in[14]), .ZN(n302) );
  INV_X1 U318 ( .A(n356), .ZN(n301) );
  INV_X1 U319 ( .A(n387), .ZN(n299) );
  OAI211_X1 U320 ( .C1(n602), .C2(n97), .A(n601), .B(n600), .ZN(a[44]) );
  AOI22_X1 U321 ( .A1(n599), .A2(n122), .B1(n128), .B2(a_in[14]), .ZN(n600) );
  INV_X1 U322 ( .A(n621), .ZN(n599) );
  AOI22_X1 U323 ( .A1(n94), .A2(n620), .B1(n625), .B2(n121), .ZN(n601) );
  INV_X1 U324 ( .A(n597), .ZN(n602) );
  OAI211_X1 U325 ( .C1(n584), .C2(n97), .A(n583), .B(n582), .ZN(a[40]) );
  AOI22_X1 U326 ( .A1(n122), .A2(n598), .B1(n128), .B2(a_in[10]), .ZN(n582) );
  AOI22_X1 U327 ( .A1(n94), .A2(n625), .B1(n597), .B2(n121), .ZN(n583) );
  OAI211_X1 U328 ( .C1(n304), .C2(n93), .A(n285), .B(n284), .ZN(neg_a[40]) );
  AOI22_X1 U329 ( .A1(n122), .A2(n283), .B1(n128), .B2(neg_a_in[10]), .ZN(n284) );
  AOI22_X1 U330 ( .A1(n94), .A2(n325), .B1(n282), .B2(n126), .ZN(n285) );
  OAI211_X1 U331 ( .C1(n588), .C2(n97), .A(n587), .B(n586), .ZN(a[41]) );
  AOI22_X1 U332 ( .A1(n122), .A2(n604), .B1(n128), .B2(a_in[11]), .ZN(n586) );
  AOI22_X1 U333 ( .A1(n94), .A2(n632), .B1(n603), .B2(n121), .ZN(n587) );
  OAI211_X1 U334 ( .C1(n310), .C2(n93), .A(n290), .B(n289), .ZN(neg_a[41]) );
  AOI22_X1 U335 ( .A1(n122), .A2(n288), .B1(n128), .B2(neg_a_in[11]), .ZN(n289) );
  AOI22_X1 U336 ( .A1(n94), .A2(n332), .B1(n287), .B2(n126), .ZN(n290) );
  OAI211_X1 U337 ( .C1(n592), .C2(n97), .A(n591), .B(n590), .ZN(a[42]) );
  AOI22_X1 U338 ( .A1(n122), .A2(n610), .B1(n128), .B2(a_in[12]), .ZN(n590) );
  AOI22_X1 U339 ( .A1(n94), .A2(n634), .B1(n611), .B2(n121), .ZN(n591) );
  OAI211_X1 U340 ( .C1(n294), .C2(n97), .A(n293), .B(n292), .ZN(neg_a[42]) );
  AOI22_X1 U341 ( .A1(n311), .A2(n122), .B1(n128), .B2(neg_a_in[12]), .ZN(n292) );
  AOI22_X1 U342 ( .A1(n94), .A2(n334), .B1(n312), .B2(n121), .ZN(n293) );
  OAI211_X1 U343 ( .C1(n298), .C2(n97), .A(n297), .B(n296), .ZN(neg_a[43]) );
  AOI22_X1 U344 ( .A1(n122), .A2(n316), .B1(n128), .B2(neg_a_in[13]), .ZN(n296) );
  AOI22_X1 U345 ( .A1(n94), .A2(n342), .B1(n317), .B2(n121), .ZN(n297) );
  OAI211_X1 U346 ( .C1(n596), .C2(n97), .A(n595), .B(n594), .ZN(a[43]) );
  AOI22_X1 U347 ( .A1(n122), .A2(n615), .B1(n128), .B2(a_in[13]), .ZN(n594) );
  AOI22_X1 U348 ( .A1(n94), .A2(n642), .B1(n616), .B2(n121), .ZN(n595) );
  OAI21_X1 U349 ( .B1(n584), .B2(n93), .A(n567), .ZN(a[36]) );
  AOI21_X1 U350 ( .B1(n94), .B2(n597), .A(n566), .ZN(n567) );
  OAI21_X1 U351 ( .B1(n565), .B2(n125), .A(n564), .ZN(n566) );
  AOI22_X1 U352 ( .A1(n122), .A2(n581), .B1(n128), .B2(a_in[6]), .ZN(n564) );
  OAI211_X1 U353 ( .C1(n304), .C2(n119), .A(n263), .B(n262), .ZN(neg_a[36]) );
  NAND2_X1 U354 ( .A1(n282), .A2(n121), .ZN(n262) );
  AOI21_X1 U355 ( .B1(n261), .B2(n126), .A(n260), .ZN(n263) );
  OAI22_X1 U356 ( .A1(n103), .A2(n259), .B1(n100), .B2(n258), .ZN(n260) );
  INV_X1 U357 ( .A(neg_a_in[34]), .ZN(n256) );
  OAI211_X1 U358 ( .C1(n298), .C2(n119), .A(n254), .B(n253), .ZN(neg_a[35]) );
  NAND2_X1 U359 ( .A1(n278), .A2(n121), .ZN(n253) );
  AOI21_X1 U360 ( .B1(n252), .B2(n126), .A(n251), .ZN(n254) );
  OAI22_X1 U361 ( .A1(n103), .A2(n250), .B1(n100), .B2(n249), .ZN(n251) );
  OAI211_X1 U362 ( .C1(n596), .C2(n119), .A(n562), .B(n561), .ZN(a[35]) );
  NAND2_X1 U363 ( .A1(n578), .A2(n121), .ZN(n561) );
  AOI21_X1 U364 ( .B1(n560), .B2(n126), .A(n559), .ZN(n562) );
  OAI22_X1 U365 ( .A1(n103), .A2(n558), .B1(n100), .B2(n557), .ZN(n559) );
  OAI211_X1 U366 ( .C1(n592), .C2(n119), .A(n553), .B(n552), .ZN(a[34]) );
  NAND2_X1 U367 ( .A1(n574), .A2(n121), .ZN(n552) );
  AOI21_X1 U368 ( .B1(n551), .B2(n126), .A(n550), .ZN(n553) );
  OAI22_X1 U369 ( .A1(n103), .A2(n549), .B1(n100), .B2(n548), .ZN(n550) );
  OAI211_X1 U370 ( .C1(n294), .C2(n91), .A(n246), .B(n245), .ZN(neg_a[34]) );
  NAND2_X1 U371 ( .A1(n274), .A2(n121), .ZN(n245) );
  AOI21_X1 U372 ( .B1(n244), .B2(n126), .A(n243), .ZN(n246) );
  OAI22_X1 U373 ( .A1(n103), .A2(n242), .B1(n100), .B2(n241), .ZN(n243) );
  OAI21_X1 U374 ( .B1(n588), .B2(n119), .A(n544), .ZN(a[33]) );
  INV_X1 U375 ( .A(n543), .ZN(n544) );
  OAI211_X1 U376 ( .C1(n542), .C2(n97), .A(n541), .B(n540), .ZN(n543) );
  AOI22_X1 U377 ( .A1(n539), .A2(n604), .B1(n122), .B2(n568), .ZN(n540) );
  AOI22_X1 U378 ( .A1(n538), .A2(n90), .B1(n128), .B2(a_in[3]), .ZN(n541) );
  OAI21_X1 U379 ( .B1(n527), .B2(n119), .A(n526), .ZN(a[31]) );
  AOI211_X1 U380 ( .C1(n126), .C2(n525), .A(n524), .B(n523), .ZN(n526) );
  OAI22_X1 U381 ( .A1(n522), .A2(n93), .B1(n100), .B2(n521), .ZN(n523) );
  NAND2_X1 U382 ( .A1(n104), .A2(n102), .ZN(n524) );
  NAND2_X1 U383 ( .A1(n539), .A2(n593), .ZN(n104) );
  INV_X1 U384 ( .A(n578), .ZN(n527) );
  OAI21_X1 U385 ( .B1(n584), .B2(n119), .A(n535), .ZN(a[32]) );
  INV_X1 U386 ( .A(n534), .ZN(n535) );
  OAI211_X1 U387 ( .C1(n533), .C2(n97), .A(n532), .B(n531), .ZN(n534) );
  AOI22_X1 U388 ( .A1(n539), .A2(n598), .B1(n122), .B2(n563), .ZN(n531) );
  AOI22_X1 U389 ( .A1(n530), .A2(n90), .B1(n128), .B2(a_in[2]), .ZN(n532) );
  INV_X1 U390 ( .A(a_in[28]), .ZN(n528) );
  OAI21_X1 U391 ( .B1(n588), .B2(n93), .A(n572), .ZN(a[37]) );
  AOI21_X1 U392 ( .B1(n94), .B2(n603), .A(n571), .ZN(n572) );
  OAI21_X1 U393 ( .B1(n570), .B2(n125), .A(n569), .ZN(n571) );
  AOI22_X1 U394 ( .A1(n122), .A2(n585), .B1(n128), .B2(a_in[7]), .ZN(n569) );
  INV_X1 U395 ( .A(a_in[29]), .ZN(n536) );
  OAI211_X1 U396 ( .C1(n310), .C2(n119), .A(n272), .B(n271), .ZN(neg_a[37]) );
  NAND2_X1 U397 ( .A1(n287), .A2(n121), .ZN(n271) );
  AOI21_X1 U398 ( .B1(n270), .B2(n126), .A(n269), .ZN(n272) );
  OAI22_X1 U399 ( .A1(n103), .A2(n268), .B1(n100), .B2(n267), .ZN(n269) );
  INV_X1 U400 ( .A(neg_a_in[35]), .ZN(n265) );
  OAI211_X1 U401 ( .C1(n592), .C2(n93), .A(n576), .B(n575), .ZN(a[38]) );
  AOI22_X1 U402 ( .A1(n122), .A2(n589), .B1(n128), .B2(a_in[8]), .ZN(n575) );
  AOI22_X1 U403 ( .A1(n94), .A2(n611), .B1(n574), .B2(n126), .ZN(n576) );
  INV_X1 U404 ( .A(a_in[30]), .ZN(n545) );
  INV_X1 U405 ( .A(a_in[32]), .ZN(n546) );
  OAI211_X1 U406 ( .C1(n294), .C2(n93), .A(n276), .B(n275), .ZN(neg_a[38]) );
  AOI22_X1 U407 ( .A1(n122), .A2(n291), .B1(n128), .B2(neg_a_in[8]), .ZN(n275)
         );
  AOI22_X1 U408 ( .A1(n94), .A2(n312), .B1(n274), .B2(n126), .ZN(n276) );
  INV_X1 U409 ( .A(neg_a_in[30]), .ZN(n239) );
  INV_X1 U410 ( .A(neg_a_in[32]), .ZN(n255) );
  OAI211_X1 U411 ( .C1(n596), .C2(n93), .A(n580), .B(n579), .ZN(a[39]) );
  AOI22_X1 U412 ( .A1(n122), .A2(n593), .B1(n128), .B2(a_in[9]), .ZN(n579) );
  AOI22_X1 U413 ( .A1(n94), .A2(n616), .B1(n578), .B2(n126), .ZN(n580) );
  INV_X1 U414 ( .A(a_in[31]), .ZN(n554) );
  INV_X1 U415 ( .A(a_in[33]), .ZN(n555) );
  OAI211_X1 U416 ( .C1(n298), .C2(n93), .A(n280), .B(n279), .ZN(neg_a[39]) );
  AOI22_X1 U417 ( .A1(n122), .A2(n295), .B1(n128), .B2(neg_a_in[9]), .ZN(n279)
         );
  AOI22_X1 U418 ( .A1(n94), .A2(n317), .B1(n278), .B2(n126), .ZN(n280) );
  INV_X1 U419 ( .A(neg_a_in[31]), .ZN(n247) );
  INV_X1 U420 ( .A(neg_a_in[33]), .ZN(n264) );
  OR2_X1 U421 ( .A1(n513), .A2(n512), .ZN(a[29]) );
  OAI22_X1 U422 ( .A1(n511), .A2(n124), .B1(n103), .B2(n537), .ZN(n512) );
  OAI22_X1 U423 ( .A1(n570), .A2(n119), .B1(n542), .B2(n93), .ZN(n513) );
  AOI21_X1 U424 ( .B1(n604), .B2(n112), .A(n538), .ZN(n570) );
  OAI211_X1 U425 ( .C1(n215), .C2(n97), .A(n214), .B(n213), .ZN(neg_a[29]) );
  NAND2_X1 U426 ( .A1(n235), .A2(n122), .ZN(n213) );
  AOI22_X1 U427 ( .A1(n270), .A2(n94), .B1(n238), .B2(n90), .ZN(n214) );
  OAI21_X1 U428 ( .B1(n134), .B2(n305), .A(n237), .ZN(n270) );
  AOI22_X1 U429 ( .A1(n498), .A2(neg_a_in[11]), .B1(neg_a_in[9]), .B2(n497), 
        .ZN(n237) );
  OAI21_X1 U430 ( .B1(n225), .B2(n91), .A(n224), .ZN(neg_a[30]) );
  AOI211_X1 U431 ( .C1(n126), .C2(n223), .A(n222), .B(n221), .ZN(n224) );
  OAI22_X1 U432 ( .A1(n220), .A2(n93), .B1(n100), .B2(n219), .ZN(n221) );
  NAND2_X1 U433 ( .A1(n105), .A2(n101), .ZN(n222) );
  NAND2_X1 U434 ( .A1(n539), .A2(n291), .ZN(n105) );
  INV_X1 U435 ( .A(n274), .ZN(n225) );
  OR2_X1 U436 ( .A1(n506), .A2(n505), .ZN(a[28]) );
  OAI22_X1 U437 ( .A1(n504), .A2(n124), .B1(n103), .B2(n529), .ZN(n505) );
  OAI22_X1 U438 ( .A1(n565), .A2(n119), .B1(n533), .B2(n93), .ZN(n506) );
  AOI21_X1 U439 ( .B1(n598), .B2(n86), .A(n530), .ZN(n565) );
  OAI211_X1 U440 ( .C1(n212), .C2(n97), .A(n211), .B(n210), .ZN(neg_a[28]) );
  NAND2_X1 U441 ( .A1(n231), .A2(n122), .ZN(n210) );
  AOI22_X1 U442 ( .A1(n261), .A2(n94), .B1(n234), .B2(n121), .ZN(n211) );
  OAI21_X1 U443 ( .B1(n134), .B2(n300), .A(n233), .ZN(n261) );
  AOI22_X1 U444 ( .A1(n498), .A2(neg_a_in[10]), .B1(neg_a_in[8]), .B2(n497), 
        .ZN(n233) );
  OAI211_X1 U445 ( .C1(n501), .C2(n97), .A(n500), .B(n499), .ZN(a[27]) );
  NAND2_X1 U446 ( .A1(n519), .A2(n122), .ZN(n499) );
  AOI22_X1 U447 ( .A1(n560), .A2(n94), .B1(n525), .B2(n121), .ZN(n500) );
  OAI21_X1 U448 ( .B1(n134), .B2(n520), .A(n522), .ZN(n560) );
  AOI22_X1 U449 ( .A1(n498), .A2(a_in[9]), .B1(n497), .B2(a_in[7]), .ZN(n522)
         );
  OAI211_X1 U450 ( .C1(n209), .C2(n97), .A(n208), .B(n207), .ZN(neg_a[27]) );
  NAND2_X1 U451 ( .A1(n226), .A2(n122), .ZN(n207) );
  AOI22_X1 U452 ( .A1(n252), .A2(n94), .B1(n230), .B2(n90), .ZN(n208) );
  OAI21_X1 U453 ( .B1(n134), .B2(n227), .A(n229), .ZN(n252) );
  AOI22_X1 U454 ( .A1(n498), .A2(neg_a_in[9]), .B1(n497), .B2(neg_a_in[7]), 
        .ZN(n229) );
  OAI211_X1 U455 ( .C1(n496), .C2(n97), .A(n495), .B(n494), .ZN(a[26]) );
  NAND2_X1 U456 ( .A1(n514), .A2(n122), .ZN(n494) );
  AOI22_X1 U457 ( .A1(n551), .A2(n94), .B1(n518), .B2(n121), .ZN(n495) );
  OAI21_X1 U458 ( .B1(n134), .B2(n515), .A(n517), .ZN(n551) );
  AOI22_X1 U459 ( .A1(n498), .A2(a_in[8]), .B1(n497), .B2(a_in[6]), .ZN(n517)
         );
  OAI211_X1 U460 ( .C1(n206), .C2(n125), .A(n205), .B(n204), .ZN(neg_a[26]) );
  NAND2_X1 U461 ( .A1(n216), .A2(n122), .ZN(n204) );
  AOI22_X1 U462 ( .A1(n244), .A2(n94), .B1(n223), .B2(n121), .ZN(n205) );
  OAI21_X1 U463 ( .B1(n134), .B2(n217), .A(n220), .ZN(n244) );
  AOI22_X1 U464 ( .A1(n498), .A2(neg_a_in[8]), .B1(n497), .B2(neg_a_in[6]), 
        .ZN(n220) );
  OAI21_X1 U465 ( .B1(n511), .B2(n93), .A(n493), .ZN(a[25]) );
  AOI211_X1 U466 ( .C1(n492), .C2(n491), .A(n490), .B(n489), .ZN(n493) );
  NOR2_X1 U467 ( .A1(n542), .A2(n119), .ZN(n489) );
  AOI21_X1 U468 ( .B1(n585), .B2(n135), .A(n488), .ZN(n542) );
  OAI22_X1 U469 ( .A1(n486), .A2(n508), .B1(n485), .B2(n509), .ZN(n490) );
  OAI211_X1 U470 ( .C1(n215), .C2(n93), .A(n203), .B(n202), .ZN(neg_a[25]) );
  NAND2_X1 U471 ( .A1(n238), .A2(n94), .ZN(n202) );
  INV_X1 U472 ( .A(n286), .ZN(n268) );
  AOI21_X1 U473 ( .B1(n235), .B2(n491), .A(n201), .ZN(n203) );
  OAI22_X1 U474 ( .A1(n486), .A2(n200), .B1(n485), .B2(n199), .ZN(n201) );
  OAI211_X1 U475 ( .C1(n501), .C2(n119), .A(n454), .B(n453), .ZN(a[19]) );
  AOI21_X1 U476 ( .B1(a_in[3]), .B2(n726), .A(n452), .ZN(n454) );
  OAI22_X1 U477 ( .A1(n487), .A2(n465), .B1(n464), .B2(n508), .ZN(n452) );
  OAI211_X1 U478 ( .C1(n209), .C2(n119), .A(n174), .B(n173), .ZN(neg_a[19]) );
  AOI21_X1 U479 ( .B1(neg_a_in[3]), .B2(n726), .A(n172), .ZN(n174) );
  OAI22_X1 U480 ( .A1(n267), .A2(n465), .B1(n464), .B2(n200), .ZN(n172) );
  OAI211_X1 U481 ( .C1(n496), .C2(n93), .A(n474), .B(n473), .ZN(a[22]) );
  NAND2_X1 U482 ( .A1(n518), .A2(n94), .ZN(n473) );
  OAI21_X1 U483 ( .B1(n549), .B2(n134), .A(n472), .ZN(n518) );
  AOI22_X1 U484 ( .A1(n498), .A2(a_in[4]), .B1(n497), .B2(a_in[2]), .ZN(n472)
         );
  INV_X1 U485 ( .A(n573), .ZN(n549) );
  AOI21_X1 U486 ( .B1(n514), .B2(n491), .A(n471), .ZN(n474) );
  OAI22_X1 U487 ( .A1(n486), .A2(n479), .B1(n485), .B2(n502), .ZN(n471) );
  OAI211_X1 U488 ( .C1(n206), .C2(n93), .A(n189), .B(n188), .ZN(neg_a[22]) );
  INV_X1 U489 ( .A(n273), .ZN(n242) );
  AOI21_X1 U490 ( .B1(n216), .B2(n491), .A(n187), .ZN(n189) );
  OAI22_X1 U491 ( .A1(n486), .A2(n258), .B1(n485), .B2(n195), .ZN(n187) );
  OAI211_X1 U492 ( .C1(n511), .C2(n119), .A(n470), .B(n469), .ZN(a[21]) );
  INV_X1 U493 ( .A(n537), .ZN(n492) );
  INV_X1 U494 ( .A(a_in[13]), .ZN(n467) );
  AOI21_X1 U495 ( .B1(a_in[5]), .B2(n726), .A(n466), .ZN(n470) );
  OAI22_X1 U496 ( .A1(n508), .A2(n465), .B1(n464), .B2(n509), .ZN(n466) );
  INV_X1 U497 ( .A(a_in[11]), .ZN(n509) );
  AOI21_X1 U498 ( .B1(n568), .B2(n135), .A(n463), .ZN(n511) );
  OAI211_X1 U499 ( .C1(n212), .C2(n119), .A(n180), .B(n179), .ZN(neg_a[20]) );
  AOI21_X1 U500 ( .B1(neg_a_in[4]), .B2(n726), .A(n178), .ZN(n180) );
  OAI22_X1 U501 ( .A1(n195), .A2(n465), .B1(n464), .B2(n194), .ZN(n178) );
  OAI211_X1 U502 ( .C1(n215), .C2(n119), .A(n186), .B(n185), .ZN(neg_a[21]) );
  AOI21_X1 U503 ( .B1(neg_a_in[5]), .B2(n726), .A(n184), .ZN(n186) );
  OAI22_X1 U504 ( .A1(n200), .A2(n465), .B1(n464), .B2(n199), .ZN(n184) );
  INV_X1 U505 ( .A(neg_a_in[11]), .ZN(n199) );
  AOI21_X1 U506 ( .B1(n183), .B2(n135), .A(n182), .ZN(n215) );
  INV_X1 U507 ( .A(n266), .ZN(n183) );
  INV_X1 U508 ( .A(neg_a_in[19]), .ZN(n327) );
  OAI211_X1 U509 ( .C1(n504), .C2(n119), .A(n461), .B(n460), .ZN(a[20]) );
  AOI21_X1 U510 ( .B1(a_in[4]), .B2(n726), .A(n457), .ZN(n461) );
  OAI22_X1 U511 ( .A1(n502), .A2(n465), .B1(n464), .B2(n503), .ZN(n457) );
  OAI211_X1 U512 ( .C1(n206), .C2(n91), .A(n169), .B(n168), .ZN(neg_a[18]) );
  AOI21_X1 U513 ( .B1(neg_a_in[2]), .B2(n726), .A(n167), .ZN(n169) );
  OAI22_X1 U514 ( .A1(n258), .A2(n465), .B1(n464), .B2(n195), .ZN(n167) );
  INV_X1 U515 ( .A(neg_a_in[6]), .ZN(n258) );
  AOI22_X1 U516 ( .A1(n166), .A2(n135), .B1(neg_a_in[0]), .B2(n498), .ZN(n206)
         );
  INV_X1 U517 ( .A(n240), .ZN(n166) );
  INV_X1 U518 ( .A(neg_a_in[14]), .ZN(n165) );
  OAI211_X1 U519 ( .C1(n496), .C2(n91), .A(n449), .B(n448), .ZN(a[18]) );
  AOI21_X1 U520 ( .B1(a_in[2]), .B2(n726), .A(n447), .ZN(n449) );
  OAI22_X1 U521 ( .A1(n479), .A2(n465), .B1(n464), .B2(n502), .ZN(n447) );
  INV_X1 U522 ( .A(n218), .ZN(n106) );
  AOI22_X1 U523 ( .A1(n446), .A2(n135), .B1(a_in[0]), .B2(n498), .ZN(n496) );
  INV_X1 U524 ( .A(n547), .ZN(n446) );
  INV_X1 U525 ( .A(a_in[16]), .ZN(n445) );
  NAND4_X1 U526 ( .A1(n164), .A2(n163), .A3(n162), .A4(n161), .ZN(neg_a[17])
         );
  AOI22_X1 U527 ( .A1(n724), .A2(neg_a_in[5]), .B1(n95), .B2(neg_a_in[7]), 
        .ZN(n162) );
  AOI22_X1 U528 ( .A1(n723), .A2(neg_a_in[13]), .B1(neg_a_in[15]), .B2(n129), 
        .ZN(n163) );
  NAND4_X1 U529 ( .A1(n444), .A2(n443), .A3(n442), .A4(n441), .ZN(a[17]) );
  AOI22_X1 U530 ( .A1(n724), .A2(a_in[5]), .B1(n95), .B2(a_in[7]), .ZN(n442)
         );
  AOI22_X1 U531 ( .A1(n723), .A2(a_in[13]), .B1(a_in[15]), .B2(n129), .ZN(n443) );
  NAND4_X1 U532 ( .A1(n434), .A2(n433), .A3(n432), .A4(n431), .ZN(a[15]) );
  NAND2_X1 U533 ( .A1(n724), .A2(a_in[3]), .ZN(n431) );
  AOI22_X1 U534 ( .A1(n92), .A2(a_in[9]), .B1(n130), .B2(a_in[13]), .ZN(n432)
         );
  AOI22_X1 U535 ( .A1(n723), .A2(a_in[11]), .B1(a_in[5]), .B2(n95), .ZN(n433)
         );
  NAND4_X1 U536 ( .A1(n160), .A2(n159), .A3(n158), .A4(n157), .ZN(neg_a[16])
         );
  AOI22_X1 U537 ( .A1(n724), .A2(neg_a_in[4]), .B1(n95), .B2(neg_a_in[6]), 
        .ZN(n158) );
  AOI22_X1 U538 ( .A1(n723), .A2(neg_a_in[12]), .B1(neg_a_in[14]), .B2(n129), 
        .ZN(n159) );
  NAND4_X1 U539 ( .A1(n438), .A2(n437), .A3(n436), .A4(n435), .ZN(a[16]) );
  AOI22_X1 U540 ( .A1(n724), .A2(a_in[4]), .B1(n95), .B2(a_in[6]), .ZN(n436)
         );
  AOI22_X1 U541 ( .A1(n723), .A2(a_in[12]), .B1(a_in[14]), .B2(n129), .ZN(n437) );
  NAND4_X1 U542 ( .A1(n156), .A2(n155), .A3(n154), .A4(n153), .ZN(neg_a[15])
         );
  NAND2_X1 U543 ( .A1(n724), .A2(neg_a_in[3]), .ZN(n153) );
  AOI22_X1 U544 ( .A1(n92), .A2(neg_a_in[9]), .B1(n129), .B2(neg_a_in[13]), 
        .ZN(n154) );
  AOI22_X1 U545 ( .A1(n723), .A2(neg_a_in[11]), .B1(neg_a_in[5]), .B2(n95), 
        .ZN(n155) );
  NAND4_X1 U546 ( .A1(n152), .A2(n151), .A3(n150), .A4(n149), .ZN(neg_a[14])
         );
  NAND2_X1 U547 ( .A1(n724), .A2(neg_a_in[2]), .ZN(n149) );
  AOI22_X1 U548 ( .A1(n92), .A2(neg_a_in[8]), .B1(n130), .B2(neg_a_in[12]), 
        .ZN(n150) );
  AOI22_X1 U549 ( .A1(n723), .A2(neg_a_in[10]), .B1(neg_a_in[4]), .B2(n95), 
        .ZN(n151) );
  NAND4_X1 U550 ( .A1(n430), .A2(n429), .A3(n428), .A4(n427), .ZN(a[14]) );
  NAND2_X1 U551 ( .A1(n724), .A2(a_in[2]), .ZN(n427) );
  AOI22_X1 U552 ( .A1(n92), .A2(a_in[8]), .B1(n130), .B2(a_in[12]), .ZN(n428)
         );
  AOI22_X1 U553 ( .A1(n723), .A2(a_in[10]), .B1(a_in[4]), .B2(n95), .ZN(n429)
         );
  AOI22_X1 U554 ( .A1(n724), .A2(a_in[1]), .B1(n95), .B2(a_in[3]), .ZN(n425)
         );
  AOI22_X1 U555 ( .A1(n92), .A2(a_in[7]), .B1(a_in[11]), .B2(n130), .ZN(n426)
         );
  AOI22_X1 U556 ( .A1(n724), .A2(neg_a_in[1]), .B1(n95), .B2(neg_a_in[3]), 
        .ZN(n147) );
  AOI22_X1 U557 ( .A1(n92), .A2(neg_a_in[7]), .B1(neg_a_in[11]), .B2(n129), 
        .ZN(n148) );
  OAI222_X1 U558 ( .A1(n236), .A2(n115), .B1(n718), .B2(n249), .C1(n228), .C2(
        n722), .ZN(neg_ax2[8]) );
  INV_X1 U559 ( .A(neg_a_in[5]), .ZN(n249) );
  OAI222_X1 U560 ( .A1(n462), .A2(n115), .B1(n718), .B2(n557), .C1(n521), .C2(
        n722), .ZN(ax2[8]) );
  INV_X1 U561 ( .A(a_in[5]), .ZN(n557) );
  NOR2_X1 U562 ( .A1(n718), .A2(n516), .ZN(a[2]) );
  NOR2_X1 U563 ( .A1(n718), .A2(n219), .ZN(neg_a[2]) );
  INV_X1 U564 ( .A(a_in[1]), .ZN(n521) );
  INV_X1 U565 ( .A(neg_a_in[1]), .ZN(n228) );
  INV_X1 U566 ( .A(neg_a_in[4]), .ZN(n241) );
  NAND2_X1 U567 ( .A1(n416), .A2(n415), .ZN(ax2[10]) );
  AOI22_X1 U568 ( .A1(n723), .A2(a_in[5]), .B1(a_in[7]), .B2(n130), .ZN(n415)
         );
  NAND2_X1 U569 ( .A1(n140), .A2(n139), .ZN(neg_ax2[10]) );
  AOI22_X1 U570 ( .A1(n723), .A2(neg_a_in[5]), .B1(neg_a_in[7]), .B2(n129), 
        .ZN(n139) );
  AOI22_X1 U571 ( .A1(n114), .A2(neg_a_in[1]), .B1(n92), .B2(neg_a_in[3]), 
        .ZN(n140) );
  OAI211_X1 U572 ( .C1(n455), .C2(n96), .A(n418), .B(n417), .ZN(ax2[11]) );
  AOI22_X1 U573 ( .A1(n723), .A2(a_in[6]), .B1(a_in[8]), .B2(n130), .ZN(n417)
         );
  AOI22_X1 U574 ( .A1(n92), .A2(a_in[4]), .B1(n95), .B2(a_in[0]), .ZN(n418) );
  OAI211_X1 U575 ( .C1(n232), .C2(n96), .A(n143), .B(n142), .ZN(neg_ax2[11])
         );
  AOI22_X1 U576 ( .A1(n723), .A2(neg_a_in[6]), .B1(neg_a_in[8]), .B2(n129), 
        .ZN(n142) );
  AOI22_X1 U577 ( .A1(n92), .A2(neg_a_in[4]), .B1(n95), .B2(neg_a_in[0]), .ZN(
        n143) );
  OAI211_X1 U578 ( .C1(n236), .C2(n96), .A(n145), .B(n144), .ZN(neg_ax2[12])
         );
  AOI22_X1 U579 ( .A1(n723), .A2(neg_a_in[7]), .B1(neg_a_in[9]), .B2(n129), 
        .ZN(n144) );
  AOI22_X1 U580 ( .A1(n92), .A2(neg_a_in[5]), .B1(n95), .B2(neg_a_in[1]), .ZN(
        n145) );
  INV_X1 U581 ( .A(neg_a_in[3]), .ZN(n236) );
  OAI211_X1 U582 ( .C1(n462), .C2(n96), .A(n420), .B(n419), .ZN(ax2[12]) );
  AOI22_X1 U583 ( .A1(n723), .A2(a_in[7]), .B1(a_in[9]), .B2(n130), .ZN(n419)
         );
  AOI22_X1 U584 ( .A1(n92), .A2(a_in[5]), .B1(n95), .B2(a_in[1]), .ZN(n420) );
  INV_X1 U585 ( .A(a_in[3]), .ZN(n462) );
  AOI22_X1 U586 ( .A1(n724), .A2(a_in[0]), .B1(n95), .B2(a_in[2]), .ZN(n422)
         );
  AOI22_X1 U587 ( .A1(n92), .A2(a_in[6]), .B1(a_in[10]), .B2(n129), .ZN(n423)
         );
  OAI21_X1 U588 ( .B1(n504), .B2(n93), .A(n484), .ZN(a[24]) );
  AOI211_X1 U589 ( .C1(n491), .C2(n483), .A(n482), .B(n481), .ZN(n484) );
  NOR2_X1 U590 ( .A1(n533), .A2(n119), .ZN(n481) );
  AOI21_X1 U591 ( .B1(n581), .B2(n86), .A(n480), .ZN(n533) );
  INV_X1 U592 ( .A(a_in[4]), .ZN(n548) );
  INV_X1 U593 ( .A(a_in[6]), .ZN(n479) );
  OAI22_X1 U594 ( .A1(n486), .A2(n502), .B1(n485), .B2(n503), .ZN(n482) );
  INV_X1 U595 ( .A(a_in[10]), .ZN(n503) );
  INV_X1 U596 ( .A(a_in[8]), .ZN(n502) );
  INV_X1 U597 ( .A(n529), .ZN(n483) );
  INV_X1 U598 ( .A(a_in[12]), .ZN(n458) );
  INV_X1 U599 ( .A(a_in[14]), .ZN(n459) );
  AOI21_X1 U600 ( .B1(n563), .B2(n135), .A(n456), .ZN(n504) );
  INV_X1 U601 ( .A(a_in[0]), .ZN(n516) );
  INV_X1 U602 ( .A(a_in[2]), .ZN(n455) );
  OAI211_X1 U603 ( .C1(n209), .C2(n93), .A(n193), .B(n192), .ZN(neg_a[23]) );
  NAND2_X1 U604 ( .A1(n230), .A2(n94), .ZN(n192) );
  NAND2_X1 U605 ( .A1(n191), .A2(n108), .ZN(n230) );
  OR2_X1 U606 ( .A1(n250), .A2(n109), .ZN(n108) );
  INV_X1 U607 ( .A(n277), .ZN(n250) );
  AOI22_X1 U608 ( .A1(n498), .A2(neg_a_in[5]), .B1(n497), .B2(neg_a_in[3]), 
        .ZN(n191) );
  AOI21_X1 U609 ( .B1(n226), .B2(n491), .A(n190), .ZN(n193) );
  OAI22_X1 U610 ( .A1(n486), .A2(n267), .B1(n485), .B2(n200), .ZN(n190) );
  INV_X1 U611 ( .A(neg_a_in[9]), .ZN(n200) );
  INV_X1 U612 ( .A(neg_a_in[7]), .ZN(n267) );
  AOI22_X1 U613 ( .A1(n171), .A2(n86), .B1(neg_a_in[1]), .B2(n498), .ZN(n209)
         );
  INV_X1 U614 ( .A(n248), .ZN(n171) );
  INV_X1 U615 ( .A(neg_a_in[15]), .ZN(n170) );
  INV_X1 U616 ( .A(neg_a_in[17]), .ZN(n181) );
  OAI211_X1 U617 ( .C1(n212), .C2(n93), .A(n198), .B(n197), .ZN(neg_a[24]) );
  NAND2_X1 U618 ( .A1(n234), .A2(n94), .ZN(n197) );
  INV_X1 U619 ( .A(n281), .ZN(n259) );
  AOI21_X1 U620 ( .B1(n231), .B2(n491), .A(n196), .ZN(n198) );
  OAI22_X1 U621 ( .A1(n486), .A2(n195), .B1(n485), .B2(n194), .ZN(n196) );
  INV_X1 U622 ( .A(neg_a_in[10]), .ZN(n194) );
  INV_X1 U623 ( .A(neg_a_in[8]), .ZN(n195) );
  AOI21_X1 U624 ( .B1(n177), .B2(n135), .A(n176), .ZN(n212) );
  INV_X1 U625 ( .A(neg_a_in[0]), .ZN(n219) );
  INV_X1 U626 ( .A(neg_a_in[2]), .ZN(n232) );
  INV_X1 U627 ( .A(n257), .ZN(n177) );
  INV_X1 U628 ( .A(neg_a_in[16]), .ZN(n175) );
  INV_X1 U629 ( .A(neg_a_in[18]), .ZN(n321) );
  OAI211_X1 U630 ( .C1(n501), .C2(n93), .A(n478), .B(n477), .ZN(a[23]) );
  NAND2_X1 U631 ( .A1(n525), .A2(n94), .ZN(n477) );
  NAND2_X1 U632 ( .A1(n476), .A2(n107), .ZN(n525) );
  OR2_X1 U633 ( .A1(n558), .A2(n109), .ZN(n107) );
  INV_X1 U634 ( .A(n577), .ZN(n558) );
  AOI22_X1 U635 ( .A1(n498), .A2(a_in[5]), .B1(n497), .B2(a_in[3]), .ZN(n476)
         );
  AOI21_X1 U636 ( .B1(n519), .B2(n491), .A(n475), .ZN(n478) );
  OAI22_X1 U637 ( .A1(n486), .A2(n487), .B1(n485), .B2(n508), .ZN(n475) );
  INV_X1 U638 ( .A(a_in[9]), .ZN(n508) );
  INV_X1 U639 ( .A(a_in[7]), .ZN(n487) );
  NOR2_X1 U640 ( .A1(n125), .A2(n109), .ZN(n491) );
  AOI22_X1 U641 ( .A1(n451), .A2(n135), .B1(a_in[1]), .B2(n498), .ZN(n501) );
  INV_X1 U642 ( .A(n556), .ZN(n451) );
  INV_X1 U643 ( .A(a_in[15]), .ZN(n468) );
  INV_X1 U644 ( .A(a_in[17]), .ZN(n450) );
  AND4_X1 U645 ( .A1(n694), .A2(n693), .A3(n692), .A4(n691), .ZN(n99) );
  INV_X1 U646 ( .A(n593), .ZN(n520) );
  INV_X1 U647 ( .A(n589), .ZN(n515) );
  INV_X1 U648 ( .A(n295), .ZN(n227) );
  INV_X1 U649 ( .A(n283), .ZN(n300) );
  INV_X1 U650 ( .A(n291), .ZN(n217) );
  INV_X1 U651 ( .A(n288), .ZN(n305) );
  OR2_X1 U652 ( .A1(n103), .A2(n240), .ZN(n101) );
  OR2_X1 U653 ( .A1(n103), .A2(n556), .ZN(n102) );
  AOI22_X1 U654 ( .A1(n92), .A2(neg_a_in[55]), .B1(n129), .B2(neg_a_in[59]), 
        .ZN(n399) );
  NAND2_X1 U655 ( .A1(n223), .A2(n605), .ZN(n188) );
  OAI222_X1 U656 ( .A1(n629), .A2(n87), .B1(n88), .B2(n733), .C1(n135), .C2(
        n628), .ZN(n661) );
  OAI222_X1 U657 ( .A1(n622), .A2(n87), .B1(n88), .B2(n732), .C1(n86), .C2(
        n621), .ZN(n655) );
  INV_X1 U658 ( .A(n371), .ZN(n397) );
  AOI211_X1 U659 ( .C1(n94), .C2(n371), .A(n354), .B(n353), .ZN(n355) );
  INV_X1 U660 ( .A(n378), .ZN(n409) );
  AOI22_X1 U661 ( .A1(n440), .A2(a_in[1]), .B1(n439), .B2(a_in[3]), .ZN(n441)
         );
  AOI22_X1 U662 ( .A1(n440), .A2(a_in[0]), .B1(n439), .B2(a_in[2]), .ZN(n435)
         );
  AOI22_X1 U663 ( .A1(n440), .A2(neg_a_in[1]), .B1(n439), .B2(neg_a_in[3]), 
        .ZN(n161) );
  AOI22_X1 U664 ( .A1(n440), .A2(neg_a_in[0]), .B1(n439), .B2(neg_a_in[2]), 
        .ZN(n157) );
  AOI22_X1 U665 ( .A1(n114), .A2(neg_a_in[6]), .B1(neg_a_in[0]), .B2(n439), 
        .ZN(n152) );
  AOI21_X1 U666 ( .B1(n661), .B2(n121), .A(n660), .ZN(n662) );
  INV_X1 U667 ( .A(n661), .ZN(n679) );
  AOI21_X1 U668 ( .B1(n655), .B2(n121), .A(n654), .ZN(n656) );
  INV_X1 U669 ( .A(n655), .ZN(n678) );
  NOR2_X1 U670 ( .A1(n718), .A2(n521), .ZN(ax2[4]) );
  AOI22_X1 U671 ( .A1(a_in[45]), .A2(n726), .B1(n725), .B2(a_in[47]), .ZN(n705) );
  AOI22_X1 U672 ( .A1(a_in[44]), .A2(n726), .B1(n725), .B2(a_in[46]), .ZN(n695) );
  AOI22_X1 U673 ( .A1(n492), .A2(n539), .B1(n725), .B2(a_in[7]), .ZN(n469) );
  AOI22_X1 U674 ( .A1(n483), .A2(n539), .B1(n725), .B2(a_in[6]), .ZN(n460) );
  AOI22_X1 U675 ( .A1(n519), .A2(n539), .B1(n725), .B2(a_in[5]), .ZN(n453) );
  AOI22_X1 U676 ( .A1(n514), .A2(n539), .B1(n725), .B2(a_in[4]), .ZN(n448) );
  AOI22_X1 U677 ( .A1(n725), .A2(neg_a_in[47]), .B1(n398), .B2(n118), .ZN(n400) );
  AOI22_X1 U678 ( .A1(n725), .A2(neg_a_in[46]), .B1(n387), .B2(n118), .ZN(n389) );
  AOI22_X1 U679 ( .A1(n235), .A2(n539), .B1(n725), .B2(neg_a_in[7]), .ZN(n185)
         );
  AOI22_X1 U680 ( .A1(n231), .A2(n539), .B1(n725), .B2(neg_a_in[6]), .ZN(n179)
         );
  AOI22_X1 U681 ( .A1(n226), .A2(n539), .B1(n725), .B2(neg_a_in[5]), .ZN(n173)
         );
  AOI22_X1 U682 ( .A1(n216), .A2(n539), .B1(n725), .B2(neg_a_in[4]), .ZN(n168)
         );
  OAI22_X1 U683 ( .A1(n510), .A2(n509), .B1(n508), .B2(n507), .ZN(n538) );
  OAI22_X1 U684 ( .A1(n510), .A2(n503), .B1(n502), .B2(n507), .ZN(n530) );
  OAI22_X1 U685 ( .A1(n510), .A2(n487), .B1(n507), .B2(n557), .ZN(n488) );
  OAI22_X1 U686 ( .A1(n510), .A2(n479), .B1(n507), .B2(n548), .ZN(n480) );
  OAI22_X1 U687 ( .A1(n510), .A2(n462), .B1(n507), .B2(n521), .ZN(n463) );
  OAI22_X1 U688 ( .A1(n510), .A2(n455), .B1(n507), .B2(n516), .ZN(n456) );
  OAI22_X1 U689 ( .A1(n510), .A2(n236), .B1(n507), .B2(n228), .ZN(n182) );
  OAI22_X1 U690 ( .A1(n510), .A2(n232), .B1(n507), .B2(n219), .ZN(n176) );
  NOR2_X1 U691 ( .A1(n141), .A2(sel[2]), .ZN(n113) );
  NAND2_X1 U692 ( .A1(n138), .A2(n137), .ZN(neg_ax2[9]) );
  AOI22_X1 U693 ( .A1(n114), .A2(neg_a_in[9]), .B1(n92), .B2(neg_a_in[11]), 
        .ZN(n164) );
  AOI22_X1 U694 ( .A1(n114), .A2(a_in[9]), .B1(n92), .B2(a_in[11]), .ZN(n444)
         );
  AOI22_X1 U695 ( .A1(n114), .A2(a_in[8]), .B1(n92), .B2(a_in[10]), .ZN(n438)
         );
  AOI22_X1 U696 ( .A1(n114), .A2(neg_a_in[8]), .B1(n92), .B2(neg_a_in[10]), 
        .ZN(n160) );
  AOI22_X1 U697 ( .A1(n114), .A2(neg_a_in[7]), .B1(neg_a_in[1]), .B2(n439), 
        .ZN(n156) );
  AOI22_X1 U698 ( .A1(n114), .A2(a_in[7]), .B1(a_in[1]), .B2(n439), .ZN(n434)
         );
  AOI22_X1 U699 ( .A1(n114), .A2(a_in[6]), .B1(a_in[0]), .B2(n439), .ZN(n430)
         );
  AOI22_X1 U700 ( .A1(n114), .A2(a_in[1]), .B1(n92), .B2(a_in[3]), .ZN(n416)
         );
  AOI22_X1 U701 ( .A1(n114), .A2(a_in[0]), .B1(n92), .B2(a_in[2]), .ZN(n414)
         );
  AOI22_X1 U702 ( .A1(n114), .A2(a_in[53]), .B1(n724), .B2(a_in[49]), .ZN(n706) );
  AOI22_X1 U703 ( .A1(n114), .A2(a_in[52]), .B1(n724), .B2(a_in[48]), .ZN(n696) );
  AOI22_X1 U704 ( .A1(n114), .A2(a_in[50]), .B1(n130), .B2(a_in[56]), .ZN(n683) );
  AOI22_X1 U705 ( .A1(a_in[5]), .A2(n114), .B1(n723), .B2(a_in[9]), .ZN(n424)
         );
  AOI22_X1 U706 ( .A1(neg_a_in[5]), .A2(n114), .B1(n723), .B2(neg_a_in[9]), 
        .ZN(n146) );
  AOI22_X1 U707 ( .A1(a_in[4]), .A2(n114), .B1(n723), .B2(a_in[8]), .ZN(n421)
         );
  AOI22_X1 U708 ( .A1(n114), .A2(neg_a_in[0]), .B1(n92), .B2(neg_a_in[2]), 
        .ZN(n138) );
  AOI22_X1 U709 ( .A1(n307), .A2(n94), .B1(n121), .B2(n332), .ZN(n309) );
  AOI22_X1 U710 ( .A1(n301), .A2(n94), .B1(n121), .B2(n325), .ZN(n303) );
  NAND2_X1 U711 ( .A1(sel[1]), .A2(sel[2]), .ZN(n218) );
  NOR2_X1 U712 ( .A1(sel[1]), .A2(sel[2]), .ZN(n605) );
  INV_X1 U713 ( .A(n723), .ZN(n117) );
  NAND2_X1 U714 ( .A1(n414), .A2(n413), .ZN(ax2[9]) );
  AOI22_X1 U715 ( .A1(n723), .A2(a_in[4]), .B1(a_in[6]), .B2(n129), .ZN(n413)
         );
  AOI22_X1 U716 ( .A1(n723), .A2(neg_a_in[4]), .B1(neg_a_in[6]), .B2(n129), 
        .ZN(n137) );
  NOR2_X1 U717 ( .A1(n87), .A2(n218), .ZN(n440) );
  NOR2_X1 U718 ( .A1(n718), .A2(n228), .ZN(neg_ax2[4]) );
  OAI211_X1 U719 ( .C1(n117), .C2(n734), .A(n653), .B(n652), .ZN(n654) );
  OAI211_X1 U720 ( .C1(n117), .C2(n736), .A(n659), .B(n658), .ZN(n660) );
  OAI211_X1 U721 ( .C1(n117), .C2(n673), .A(n672), .B(n671), .ZN(n674) );
  OAI211_X1 U722 ( .C1(n117), .C2(n392), .A(n374), .B(n373), .ZN(n375) );
  OAI211_X1 U723 ( .C1(n117), .C2(n404), .A(n381), .B(n380), .ZN(n382) );
  OAI211_X1 U724 ( .C1(n117), .C2(n728), .A(n360), .B(n359), .ZN(n361) );
  OAI211_X1 U725 ( .C1(n117), .C2(n730), .A(n366), .B(n365), .ZN(n367) );
  OAI211_X1 U726 ( .C1(n117), .C2(n666), .A(n665), .B(n664), .ZN(n667) );
  OAI22_X1 U727 ( .A1(n718), .A2(n462), .B1(n115), .B2(n521), .ZN(ax2[6]) );
  OAI222_X1 U728 ( .A1(n722), .A2(n219), .B1(n718), .B2(n241), .C1(n232), .C2(
        n116), .ZN(neg_ax2[7]) );
  OAI22_X1 U729 ( .A1(n718), .A2(n455), .B1(n116), .B2(n516), .ZN(ax2[5]) );
  OAI22_X1 U730 ( .A1(n718), .A2(n236), .B1(n115), .B2(n228), .ZN(neg_ax2[6])
         );
  OAI222_X1 U731 ( .A1(n722), .A2(n516), .B1(n718), .B2(n548), .C1(n455), .C2(
        n116), .ZN(ax2[7]) );
  OAI22_X1 U732 ( .A1(n718), .A2(n232), .B1(n219), .B2(n116), .ZN(neg_ax2[5])
         );
  AOI222_X1 U733 ( .A1(neg_a_in[47]), .A2(n329), .B1(neg_a_in[45]), .B2(n98), 
        .C1(n134), .C2(n328), .ZN(n379) );
  AOI222_X1 U734 ( .A1(neg_a_in[46]), .A2(n329), .B1(n98), .B2(neg_a_in[44]), 
        .C1(n134), .C2(n322), .ZN(n372) );
  OAI222_X1 U735 ( .A1(n350), .A2(n112), .B1(n87), .B2(n727), .C1(n88), .C2(
        n728), .ZN(n371) );
  OAI222_X1 U736 ( .A1(n357), .A2(n112), .B1(n87), .B2(n729), .C1(n88), .C2(
        n730), .ZN(n378) );
  OAI22_X1 U737 ( .A1(n87), .A2(n733), .B1(n88), .B2(n736), .ZN(n645) );
  OAI22_X1 U738 ( .A1(n87), .A2(n731), .B1(n88), .B2(n727), .ZN(n335) );
  OAI22_X1 U739 ( .A1(n87), .A2(n735), .B1(n88), .B2(n729), .ZN(n343) );
  OAI22_X1 U740 ( .A1(n87), .A2(n732), .B1(n88), .B2(n734), .ZN(n635) );
  NOR2_X1 U741 ( .A1(n88), .A2(n218), .ZN(n439) );
  INV_X1 U742 ( .A(n643), .ZN(n329) );
  INV_X1 U743 ( .A(n605), .ZN(n120) );
  INV_X1 U744 ( .A(n103), .ZN(n123) );
  NAND3_X1 U745 ( .A1(n148), .A2(n147), .A3(n146), .ZN(neg_a[13]) );
  MUX2_X1 U746 ( .A(n175), .B(n165), .S(n132), .Z(n240) );
  MUX2_X1 U747 ( .A(neg_a_in[12]), .B(neg_a_in[10]), .S(n132), .Z(n216) );
  MUX2_X1 U748 ( .A(n181), .B(n170), .S(n132), .Z(n248) );
  MUX2_X1 U749 ( .A(neg_a_in[13]), .B(neg_a_in[11]), .S(n111), .Z(n226) );
  MUX2_X1 U750 ( .A(n321), .B(n175), .S(n132), .Z(n257) );
  MUX2_X1 U751 ( .A(neg_a_in[14]), .B(neg_a_in[12]), .S(n132), .Z(n231) );
  MUX2_X1 U752 ( .A(n327), .B(n181), .S(n132), .Z(n266) );
  MUX2_X1 U753 ( .A(neg_a_in[15]), .B(neg_a_in[13]), .S(n132), .Z(n235) );
  MUX2_X1 U754 ( .A(neg_a_in[20]), .B(neg_a_in[18]), .S(n111), .Z(n273) );
  MUX2_X1 U755 ( .A(neg_a_in[21]), .B(neg_a_in[19]), .S(n132), .Z(n277) );
  MUX2_X1 U756 ( .A(neg_a_in[22]), .B(neg_a_in[20]), .S(n111), .Z(n281) );
  MUX2_X1 U757 ( .A(neg_a_in[23]), .B(neg_a_in[21]), .S(n111), .Z(n286) );
  MUX2_X1 U758 ( .A(neg_a_in[24]), .B(neg_a_in[22]), .S(n132), .Z(n291) );
  MUX2_X1 U759 ( .A(neg_a_in[25]), .B(neg_a_in[23]), .S(n132), .Z(n295) );
  MUX2_X1 U760 ( .A(neg_a_in[26]), .B(neg_a_in[24]), .S(n132), .Z(n283) );
  MUX2_X1 U761 ( .A(neg_a_in[27]), .B(neg_a_in[25]), .S(n132), .Z(n288) );
  MUX2_X1 U762 ( .A(neg_a_in[28]), .B(neg_a_in[26]), .S(n111), .Z(n311) );
  MUX2_X1 U763 ( .A(n216), .B(n311), .S(n135), .Z(n274) );
  MUX2_X1 U764 ( .A(neg_a_in[29]), .B(neg_a_in[27]), .S(n111), .Z(n316) );
  MUX2_X1 U765 ( .A(n226), .B(n316), .S(n112), .Z(n278) );
  MUX2_X1 U766 ( .A(neg_a_in[30]), .B(neg_a_in[28]), .S(n111), .Z(n322) );
  MUX2_X1 U767 ( .A(n231), .B(n322), .S(n112), .Z(n282) );
  MUX2_X1 U768 ( .A(neg_a_in[31]), .B(neg_a_in[29]), .S(n132), .Z(n328) );
  MUX2_X1 U769 ( .A(n235), .B(n328), .S(n86), .Z(n287) );
  MUX2_X1 U770 ( .A(n255), .B(n239), .S(n111), .Z(n313) );
  MUX2_X1 U771 ( .A(n313), .B(n240), .S(n134), .Z(n294) );
  MUX2_X1 U772 ( .A(n264), .B(n247), .S(n132), .Z(n318) );
  MUX2_X1 U773 ( .A(n318), .B(n248), .S(n134), .Z(n298) );
  MUX2_X1 U774 ( .A(n256), .B(n255), .S(n89), .Z(n350) );
  MUX2_X1 U775 ( .A(n350), .B(n257), .S(n134), .Z(n304) );
  MUX2_X1 U776 ( .A(n265), .B(n264), .S(n132), .Z(n357) );
  MUX2_X1 U777 ( .A(n357), .B(n266), .S(n134), .Z(n310) );
  MUX2_X1 U778 ( .A(neg_a_in[36]), .B(neg_a_in[34]), .S(n132), .Z(n411) );
  MUX2_X1 U779 ( .A(n411), .B(n273), .S(n134), .Z(n312) );
  MUX2_X1 U780 ( .A(neg_a_in[37]), .B(neg_a_in[35]), .S(n132), .Z(n713) );
  MUX2_X1 U781 ( .A(n713), .B(n277), .S(n134), .Z(n317) );
  MUX2_X1 U782 ( .A(neg_a_in[38]), .B(neg_a_in[36]), .S(n131), .Z(n395) );
  MUX2_X1 U783 ( .A(n395), .B(n281), .S(n134), .Z(n325) );
  MUX2_X1 U784 ( .A(neg_a_in[39]), .B(neg_a_in[37]), .S(n111), .Z(n407) );
  MUX2_X1 U785 ( .A(n407), .B(n286), .S(n134), .Z(n332) );
  MUX2_X1 U786 ( .A(neg_a_in[40]), .B(neg_a_in[38]), .S(n131), .Z(n412) );
  MUX2_X1 U787 ( .A(n412), .B(n291), .S(n134), .Z(n334) );
  MUX2_X1 U788 ( .A(neg_a_in[41]), .B(neg_a_in[39]), .S(n111), .Z(n714) );
  MUX2_X1 U789 ( .A(n714), .B(n295), .S(n134), .Z(n342) );
  MUX2_X1 U790 ( .A(neg_a_in[42]), .B(neg_a_in[40]), .S(n131), .Z(n387) );
  MUX2_X1 U791 ( .A(n300), .B(n299), .S(n112), .Z(n356) );
  MUX2_X1 U792 ( .A(neg_a_in[43]), .B(neg_a_in[41]), .S(n132), .Z(n398) );
  MUX2_X1 U793 ( .A(n306), .B(n305), .S(n134), .Z(n358) );
  MUX2_X1 U794 ( .A(neg_a_in[44]), .B(neg_a_in[42]), .S(n131), .Z(n410) );
  MUX2_X1 U795 ( .A(n410), .B(n311), .S(n134), .Z(n339) );
  MUX2_X1 U796 ( .A(neg_a_in[45]), .B(neg_a_in[43]), .S(n131), .Z(n712) );
  MUX2_X1 U797 ( .A(n712), .B(n316), .S(n134), .Z(n347) );
  NAND3_X1 U798 ( .A1(n423), .A2(n422), .A3(n421), .ZN(a[12]) );
  NAND3_X1 U799 ( .A1(n426), .A2(n425), .A3(n424), .ZN(a[13]) );
  MUX2_X1 U800 ( .A(n445), .B(n459), .S(n132), .Z(n547) );
  MUX2_X1 U801 ( .A(a_in[12]), .B(a_in[10]), .S(n132), .Z(n514) );
  MUX2_X1 U802 ( .A(n450), .B(n468), .S(n132), .Z(n556) );
  MUX2_X1 U803 ( .A(a_in[13]), .B(a_in[11]), .S(n111), .Z(n519) );
  MUX2_X1 U804 ( .A(a_in[18]), .B(a_in[16]), .S(n132), .Z(n563) );
  MUX2_X1 U805 ( .A(n459), .B(n458), .S(n132), .Z(n529) );
  MUX2_X1 U806 ( .A(a_in[19]), .B(a_in[17]), .S(n132), .Z(n568) );
  MUX2_X1 U807 ( .A(n468), .B(n467), .S(n132), .Z(n537) );
  MUX2_X1 U808 ( .A(a_in[20]), .B(a_in[18]), .S(n132), .Z(n573) );
  MUX2_X1 U809 ( .A(a_in[21]), .B(a_in[19]), .S(n132), .Z(n577) );
  MUX2_X1 U810 ( .A(a_in[22]), .B(a_in[20]), .S(n132), .Z(n581) );
  MUX2_X1 U811 ( .A(a_in[23]), .B(a_in[21]), .S(n111), .Z(n585) );
  MUX2_X1 U812 ( .A(a_in[24]), .B(a_in[22]), .S(n131), .Z(n589) );
  MUX2_X1 U813 ( .A(a_in[25]), .B(a_in[23]), .S(n111), .Z(n593) );
  MUX2_X1 U814 ( .A(a_in[26]), .B(a_in[24]), .S(n132), .Z(n598) );
  MUX2_X1 U815 ( .A(a_in[27]), .B(a_in[25]), .S(n132), .Z(n604) );
  MUX2_X1 U816 ( .A(a_in[28]), .B(a_in[26]), .S(n131), .Z(n610) );
  MUX2_X1 U817 ( .A(n514), .B(n610), .S(n112), .Z(n574) );
  MUX2_X1 U818 ( .A(a_in[29]), .B(a_in[27]), .S(n111), .Z(n615) );
  MUX2_X1 U819 ( .A(n519), .B(n615), .S(n112), .Z(n578) );
  MUX2_X1 U820 ( .A(n545), .B(n528), .S(n132), .Z(n621) );
  MUX2_X1 U821 ( .A(n529), .B(n621), .S(n86), .Z(n584) );
  MUX2_X1 U822 ( .A(n554), .B(n536), .S(n132), .Z(n628) );
  MUX2_X1 U823 ( .A(n628), .B(n537), .S(n134), .Z(n588) );
  MUX2_X1 U824 ( .A(n546), .B(n545), .S(n131), .Z(n612) );
  MUX2_X1 U825 ( .A(n612), .B(n547), .S(n134), .Z(n592) );
  MUX2_X1 U826 ( .A(n555), .B(n554), .S(n131), .Z(n617) );
  MUX2_X1 U827 ( .A(n617), .B(n556), .S(n134), .Z(n596) );
  MUX2_X1 U828 ( .A(a_in[34]), .B(a_in[32]), .S(n132), .Z(n690) );
  MUX2_X1 U829 ( .A(n690), .B(n563), .S(n134), .Z(n597) );
  MUX2_X1 U830 ( .A(a_in[35]), .B(a_in[33]), .S(n111), .Z(n700) );
  MUX2_X1 U831 ( .A(n700), .B(n568), .S(n134), .Z(n603) );
  MUX2_X1 U832 ( .A(a_in[36]), .B(a_in[34]), .S(n132), .Z(n711) );
  MUX2_X1 U833 ( .A(n711), .B(n573), .S(n134), .Z(n611) );
  MUX2_X1 U834 ( .A(a_in[37]), .B(a_in[35]), .S(n132), .Z(n720) );
  MUX2_X1 U835 ( .A(n720), .B(n577), .S(n134), .Z(n616) );
  MUX2_X1 U836 ( .A(a_in[38]), .B(a_in[36]), .S(n89), .Z(n689) );
  MUX2_X1 U837 ( .A(n689), .B(n581), .S(n134), .Z(n625) );
  MUX2_X1 U838 ( .A(a_in[39]), .B(a_in[37]), .S(n132), .Z(n699) );
  MUX2_X1 U839 ( .A(n699), .B(n585), .S(n134), .Z(n632) );
  MUX2_X1 U840 ( .A(a_in[40]), .B(a_in[38]), .S(n132), .Z(n710) );
  MUX2_X1 U841 ( .A(n710), .B(n589), .S(n134), .Z(n634) );
  MUX2_X1 U842 ( .A(a_in[41]), .B(a_in[39]), .S(n89), .Z(n716) );
  MUX2_X1 U843 ( .A(n716), .B(n593), .S(n134), .Z(n642) );
  MUX2_X1 U844 ( .A(a_in[42]), .B(a_in[40]), .S(n89), .Z(n688) );
  MUX2_X1 U845 ( .A(n598), .B(n688), .S(n112), .Z(n620) );
  MUX2_X1 U846 ( .A(a_in[43]), .B(a_in[41]), .S(n132), .Z(n698) );
  MUX2_X1 U847 ( .A(n604), .B(n698), .S(n112), .Z(n627) );
  MUX2_X1 U848 ( .A(a_in[44]), .B(a_in[42]), .S(n131), .Z(n709) );
  MUX2_X1 U849 ( .A(n709), .B(n610), .S(n134), .Z(n639) );
  MUX2_X1 U850 ( .A(a_in[45]), .B(a_in[43]), .S(n132), .Z(n715) );
  MUX2_X1 U851 ( .A(n715), .B(n615), .S(n134), .Z(n649) );
  INV_X1 U852 ( .A(neg_a_in[46]), .ZN(n731) );
  INV_X1 U853 ( .A(neg_a_in[47]), .ZN(n735) );
  INV_X1 U854 ( .A(neg_a_in[48]), .ZN(n727) );
  INV_X1 U855 ( .A(neg_a_in[49]), .ZN(n729) );
  INV_X1 U856 ( .A(neg_a_in[50]), .ZN(n728) );
  INV_X1 U857 ( .A(neg_a_in[51]), .ZN(n730) );
  INV_X1 U858 ( .A(a_in[46]), .ZN(n732) );
  INV_X1 U859 ( .A(a_in[47]), .ZN(n733) );
  INV_X1 U860 ( .A(a_in[48]), .ZN(n734) );
  INV_X1 U861 ( .A(a_in[49]), .ZN(n736) );
endmodule


module dlx_syn ( clk, rst, btb_cache_update_line, btb_cache_update_data, 
        btb_cache_hit_read, btb_cache_hit_rw, btb_cache_read_address, 
        btb_cache_rw_address, btb_cache_data_in, btb_cache_data_out_read, 
        btb_cache_data_out_rw, pc_out, instr_if, dcache_hit, dcache_update, 
        dcache_update_type, dcache_data_in, dcache_address, dcache_data_out, 
        ram_update, ram_to_cache_data, cache_to_ram_data, cpu_cache_address, 
        evicted_cache_address, ram_rw, ram_address, ram_data_in, ram_data_out, 
        pc_en, predicted_taken, taken, wp_en, hilo_wr_en, rd, wp_data, 
        wp_alu_data_high );
  output [29:0] btb_cache_read_address;
  output [29:0] btb_cache_rw_address;
  output [31:0] btb_cache_data_in;
  input [31:0] btb_cache_data_out_read;
  input [31:0] btb_cache_data_out_rw;
  output [29:0] pc_out;
  input [31:0] instr_if;
  output [1:0] dcache_update_type;
  input [31:0] dcache_data_in;
  output [31:0] dcache_address;
  output [31:0] dcache_data_out;
  output [31:0] ram_to_cache_data;
  input [31:0] cache_to_ram_data;
  input [31:0] cpu_cache_address;
  input [31:0] evicted_cache_address;
  output [7:0] ram_address;
  output [31:0] ram_data_in;
  input [31:0] ram_data_out;
  output [4:0] rd;
  output [31:0] wp_data;
  output [31:0] wp_alu_data_high;
  input clk, rst, btb_cache_hit_read, btb_cache_hit_rw, dcache_hit, ram_update;
  output btb_cache_update_line, btb_cache_update_data, dcache_update, ram_rw,
         pc_en, predicted_taken, taken, wp_en, hilo_wr_en;
  wire   n7533, n7534, n7535, n7536, n7537, n7538, btb_addr_known_if,
         j_instr_id, is_signed_id, sign_ext_sel_id, b_selector_id,
         data_tbs_selector_id, sub_add_exe, op_sign_exe, en_b_exe,
         rst_exe_mem_regs, ld_sign_mem, alu_data_tbs_selector, en_alu_mem,
         en_cache_mem, rst_mem_wb_regs, cpu_is_reading, wr_mem,
         \dp/cache_data_mem_wb_int[31] , \dp/cache_data_mem_wb_int[30] ,
         \dp/cache_data_mem_wb_int[29] , \dp/cache_data_mem_wb_int[28] ,
         \dp/cache_data_mem_wb_int[27] , \dp/cache_data_mem_wb_int[26] ,
         \dp/cache_data_mem_wb_int[25] , \dp/cache_data_mem_wb_int[24] ,
         \dp/cache_data_mem_wb_int[23] , \dp/cache_data_mem_wb_int[22] ,
         \dp/cache_data_mem_wb_int[21] , \dp/cache_data_mem_wb_int[20] ,
         \dp/cache_data_mem_wb_int[19] , \dp/cache_data_mem_wb_int[18] ,
         \dp/cache_data_mem_wb_int[17] , \dp/cache_data_mem_wb_int[16] ,
         \dp/cache_data_mem_wb_int[15] , \dp/cache_data_mem_wb_int[14] ,
         \dp/cache_data_mem_wb_int[13] , \dp/cache_data_mem_wb_int[12] ,
         \dp/cache_data_mem_wb_int[11] , \dp/cache_data_mem_wb_int[10] ,
         \dp/cache_data_mem_wb_int[9] , \dp/cache_data_mem_wb_int[8] ,
         \dp/cache_data_mem_wb_int[7] , \dp/cache_data_mem_wb_int[6] ,
         \dp/cache_data_mem_wb_int[5] , \dp/cache_data_mem_wb_int[4] ,
         \dp/cache_data_mem_wb_int[3] , \dp/cache_data_mem_wb_int[2] ,
         \dp/cache_data_mem_wb_int[1] , \dp/cache_data_mem_wb_int[0] ,
         \dp/cache_in_mem_int[7] , \dp/cache_in_mem_int[6] ,
         \dp/cache_in_mem_int[5] , \dp/cache_in_mem_int[4] ,
         \dp/cache_in_mem_int[3] , \dp/cache_in_mem_int[2] ,
         \dp/cache_in_mem_int[1] , \dp/cache_in_mem_int[0] ,
         \dp/mul_feedback_exe_mem_int[62] , \dp/mul_feedback_exe_mem_int[61] ,
         \dp/mul_feedback_exe_mem_int[60] , \dp/mul_feedback_exe_mem_int[59] ,
         \dp/mul_feedback_exe_mem_int[58] , \dp/mul_feedback_exe_mem_int[57] ,
         \dp/mul_feedback_exe_mem_int[56] , \dp/mul_feedback_exe_mem_int[55] ,
         \dp/mul_feedback_exe_mem_int[54] , \dp/mul_feedback_exe_mem_int[53] ,
         \dp/mul_feedback_exe_mem_int[52] , \dp/mul_feedback_exe_mem_int[51] ,
         \dp/mul_feedback_exe_mem_int[50] , \dp/mul_feedback_exe_mem_int[49] ,
         \dp/mul_feedback_exe_mem_int[48] , \dp/mul_feedback_exe_mem_int[47] ,
         \dp/mul_feedback_exe_mem_int[46] , \dp/mul_feedback_exe_mem_int[45] ,
         \dp/mul_feedback_exe_mem_int[44] , \dp/mul_feedback_exe_mem_int[43] ,
         \dp/mul_feedback_exe_mem_int[42] , \dp/mul_feedback_exe_mem_int[41] ,
         \dp/mul_feedback_exe_mem_int[40] , \dp/mul_feedback_exe_mem_int[39] ,
         \dp/mul_feedback_exe_mem_int[38] , \dp/mul_feedback_exe_mem_int[37] ,
         \dp/mul_feedback_exe_mem_int[36] , \dp/mul_feedback_exe_mem_int[35] ,
         \dp/mul_feedback_exe_mem_int[34] , \dp/mul_feedback_exe_mem_int[33] ,
         \dp/mul_feedback_exe_mem_int[32] , \dp/mul_feedback_exe_mem_int[31] ,
         \dp/mul_feedback_exe_mem_int[30] , \dp/mul_feedback_exe_mem_int[29] ,
         \dp/mul_feedback_exe_mem_int[28] , \dp/mul_feedback_exe_mem_int[27] ,
         \dp/mul_feedback_exe_mem_int[26] , \dp/mul_feedback_exe_mem_int[25] ,
         \dp/mul_feedback_exe_mem_int[24] , \dp/mul_feedback_exe_mem_int[23] ,
         \dp/mul_feedback_exe_mem_int[22] , \dp/mul_feedback_exe_mem_int[21] ,
         \dp/mul_feedback_exe_mem_int[20] , \dp/mul_feedback_exe_mem_int[19] ,
         \dp/mul_feedback_exe_mem_int[18] , \dp/mul_feedback_exe_mem_int[17] ,
         \dp/mul_feedback_exe_mem_int[16] , \dp/mul_feedback_exe_mem_int[15] ,
         \dp/mul_feedback_exe_mem_int[14] , \dp/mul_feedback_exe_mem_int[13] ,
         \dp/mul_feedback_exe_mem_int[12] , \dp/mul_feedback_exe_mem_int[11] ,
         \dp/mul_feedback_exe_mem_int[10] , \dp/mul_feedback_exe_mem_int[9] ,
         \dp/mul_feedback_exe_mem_int[8] , \dp/mul_feedback_exe_mem_int[7] ,
         \dp/mul_feedback_exe_mem_int[6] , \dp/mul_feedback_exe_mem_int[5] ,
         \dp/mul_feedback_exe_mem_int[4] , \dp/mul_feedback_exe_mem_int[3] ,
         \dp/mul_feedback_exe_mem_int[2] , \dp/mul_feedback_exe_mem_int[1] ,
         \dp/mul_feedback_exe_mem_int[0] , \dp/b10_1_mult_id_exe_int[1] ,
         \dp/b_mult_id_exe_int[2] , \dp/a_neg_mult_id_exe_int[63] ,
         \dp/a_neg_mult_id_exe_int[62] , \dp/a_neg_mult_id_exe_int[61] ,
         \dp/a_neg_mult_id_exe_int[60] , \dp/a_neg_mult_id_exe_int[59] ,
         \dp/a_neg_mult_id_exe_int[58] , \dp/a_neg_mult_id_exe_int[57] ,
         \dp/a_neg_mult_id_exe_int[56] , \dp/a_neg_mult_id_exe_int[55] ,
         \dp/a_neg_mult_id_exe_int[54] , \dp/a_neg_mult_id_exe_int[53] ,
         \dp/a_neg_mult_id_exe_int[52] , \dp/a_neg_mult_id_exe_int[51] ,
         \dp/a_neg_mult_id_exe_int[50] , \dp/a_neg_mult_id_exe_int[49] ,
         \dp/a_neg_mult_id_exe_int[48] , \dp/a_neg_mult_id_exe_int[47] ,
         \dp/a_neg_mult_id_exe_int[46] , \dp/a_neg_mult_id_exe_int[45] ,
         \dp/a_neg_mult_id_exe_int[44] , \dp/a_neg_mult_id_exe_int[43] ,
         \dp/a_neg_mult_id_exe_int[42] , \dp/a_neg_mult_id_exe_int[41] ,
         \dp/a_neg_mult_id_exe_int[40] , \dp/a_neg_mult_id_exe_int[39] ,
         \dp/a_neg_mult_id_exe_int[38] , \dp/a_neg_mult_id_exe_int[37] ,
         \dp/a_neg_mult_id_exe_int[36] , \dp/a_neg_mult_id_exe_int[35] ,
         \dp/a_neg_mult_id_exe_int[34] , \dp/a_neg_mult_id_exe_int[33] ,
         \dp/a_neg_mult_id_exe_int[32] , \dp/a_neg_mult_id_exe_int[31] ,
         \dp/a_neg_mult_id_exe_int[30] , \dp/a_neg_mult_id_exe_int[29] ,
         \dp/a_neg_mult_id_exe_int[28] , \dp/a_neg_mult_id_exe_int[27] ,
         \dp/a_neg_mult_id_exe_int[26] , \dp/a_neg_mult_id_exe_int[25] ,
         \dp/a_neg_mult_id_exe_int[24] , \dp/a_neg_mult_id_exe_int[23] ,
         \dp/a_neg_mult_id_exe_int[22] , \dp/a_neg_mult_id_exe_int[21] ,
         \dp/a_neg_mult_id_exe_int[20] , \dp/a_neg_mult_id_exe_int[19] ,
         \dp/a_neg_mult_id_exe_int[18] , \dp/a_neg_mult_id_exe_int[17] ,
         \dp/a_neg_mult_id_exe_int[16] , \dp/a_neg_mult_id_exe_int[15] ,
         \dp/a_neg_mult_id_exe_int[14] , \dp/a_neg_mult_id_exe_int[13] ,
         \dp/a_neg_mult_id_exe_int[12] , \dp/a_neg_mult_id_exe_int[11] ,
         \dp/a_neg_mult_id_exe_int[10] , \dp/a_neg_mult_id_exe_int[9] ,
         \dp/a_neg_mult_id_exe_int[8] , \dp/a_neg_mult_id_exe_int[7] ,
         \dp/a_neg_mult_id_exe_int[6] , \dp/a_neg_mult_id_exe_int[5] ,
         \dp/a_neg_mult_id_exe_int[4] , \dp/a_neg_mult_id_exe_int[3] ,
         \dp/a_neg_mult_id_exe_int[2] , \dp/a_neg_mult_id_exe_int[1] ,
         \dp/a_neg_mult_id_exe_int[0] , \dp/a_mult_id_exe_int[63] ,
         \dp/a_mult_id_exe_int[62] , \dp/a_mult_id_exe_int[61] ,
         \dp/a_mult_id_exe_int[60] , \dp/a_mult_id_exe_int[59] ,
         \dp/a_mult_id_exe_int[58] , \dp/a_mult_id_exe_int[57] ,
         \dp/a_mult_id_exe_int[56] , \dp/a_mult_id_exe_int[55] ,
         \dp/a_mult_id_exe_int[54] , \dp/a_mult_id_exe_int[53] ,
         \dp/a_mult_id_exe_int[52] , \dp/a_mult_id_exe_int[51] ,
         \dp/a_mult_id_exe_int[50] , \dp/a_mult_id_exe_int[49] ,
         \dp/a_mult_id_exe_int[48] , \dp/a_mult_id_exe_int[47] ,
         \dp/a_mult_id_exe_int[46] , \dp/a_mult_id_exe_int[45] ,
         \dp/a_mult_id_exe_int[44] , \dp/a_mult_id_exe_int[43] ,
         \dp/a_mult_id_exe_int[42] , \dp/a_mult_id_exe_int[41] ,
         \dp/a_mult_id_exe_int[40] , \dp/a_mult_id_exe_int[39] ,
         \dp/a_mult_id_exe_int[38] , \dp/a_mult_id_exe_int[37] ,
         \dp/a_mult_id_exe_int[36] , \dp/a_mult_id_exe_int[35] ,
         \dp/a_mult_id_exe_int[34] , \dp/a_mult_id_exe_int[33] ,
         \dp/a_mult_id_exe_int[32] , \dp/a_mult_id_exe_int[31] ,
         \dp/a_mult_id_exe_int[30] , \dp/a_mult_id_exe_int[29] ,
         \dp/a_mult_id_exe_int[28] , \dp/a_mult_id_exe_int[27] ,
         \dp/a_mult_id_exe_int[26] , \dp/a_mult_id_exe_int[25] ,
         \dp/a_mult_id_exe_int[24] , \dp/a_mult_id_exe_int[23] ,
         \dp/a_mult_id_exe_int[22] , \dp/a_mult_id_exe_int[21] ,
         \dp/a_mult_id_exe_int[20] , \dp/a_mult_id_exe_int[19] ,
         \dp/a_mult_id_exe_int[18] , \dp/a_mult_id_exe_int[17] ,
         \dp/a_mult_id_exe_int[16] , \dp/a_mult_id_exe_int[15] ,
         \dp/a_mult_id_exe_int[14] , \dp/a_mult_id_exe_int[13] ,
         \dp/a_mult_id_exe_int[12] , \dp/a_mult_id_exe_int[11] ,
         \dp/a_mult_id_exe_int[10] , \dp/a_mult_id_exe_int[9] ,
         \dp/a_mult_id_exe_int[8] , \dp/a_mult_id_exe_int[7] ,
         \dp/a_mult_id_exe_int[6] , \dp/a_mult_id_exe_int[5] ,
         \dp/a_mult_id_exe_int[4] , \dp/a_mult_id_exe_int[3] ,
         \dp/a_mult_id_exe_int[2] , \dp/a_mult_id_exe_int[1] ,
         \dp/a_mult_id_exe_int[0] , \dp/b_adder_id_exe_int[31] ,
         \dp/b_adder_id_exe_int[25] , \dp/b_adder_id_exe_int[24] ,
         \dp/b_adder_id_exe_int[23] , \dp/b_adder_id_exe_int[22] ,
         \dp/b_adder_id_exe_int[21] , \dp/b_adder_id_exe_int[20] ,
         \dp/b_adder_id_exe_int[19] , \dp/b_adder_id_exe_int[18] ,
         \dp/b_adder_id_exe_int[17] , \dp/b_adder_id_exe_int[16] ,
         \dp/b_adder_id_exe_int[15] , \dp/b_adder_id_exe_int[14] ,
         \dp/b_adder_id_exe_int[13] , \dp/b_adder_id_exe_int[12] ,
         \dp/b_adder_id_exe_int[11] , \dp/b_adder_id_exe_int[10] ,
         \dp/b_adder_id_exe_int[9] , \dp/b_adder_id_exe_int[8] ,
         \dp/b_adder_id_exe_int[7] , \dp/b_adder_id_exe_int[6] ,
         \dp/b_adder_id_exe_int[5] , \dp/b_adder_id_exe_int[4] ,
         \dp/b_adder_id_exe_int[3] , \dp/b_adder_id_exe_int[2] ,
         \dp/b_adder_id_exe_int[1] , \dp/b_adder_id_exe_int[0] ,
         \dp/imm_id_exe_int[31] , \dp/imm_id_exe_int[30] ,
         \dp/imm_id_exe_int[24] , \dp/imm_id_exe_int[23] ,
         \dp/imm_id_exe_int[22] , \dp/imm_id_exe_int[21] ,
         \dp/imm_id_exe_int[16] , \dp/imm_id_exe_int[15] ,
         \dp/imm_id_exe_int[8] , \dp/imm_id_exe_int[6] ,
         \dp/imm_id_exe_int[4] , \dp/imm_id_exe_int[2] ,
         \dp/op_b_id_ex_int[31] , \dp/op_b_id_ex_int[30] ,
         \dp/op_b_id_ex_int[29] , \dp/op_b_id_ex_int[28] ,
         \dp/op_b_id_ex_int[27] , \dp/op_b_id_ex_int[26] ,
         \dp/op_b_id_ex_int[25] , \dp/op_b_id_ex_int[24] ,
         \dp/op_b_id_ex_int[23] , \dp/op_b_id_ex_int[22] ,
         \dp/op_b_id_ex_int[21] , \dp/op_b_id_ex_int[20] ,
         \dp/op_b_id_ex_int[19] , \dp/op_b_id_ex_int[18] ,
         \dp/op_b_id_ex_int[17] , \dp/op_b_id_ex_int[16] ,
         \dp/op_b_id_ex_int[15] , \dp/op_b_id_ex_int[14] ,
         \dp/op_b_id_ex_int[13] , \dp/op_b_id_ex_int[12] ,
         \dp/op_b_id_ex_int[11] , \dp/op_b_id_ex_int[10] ,
         \dp/op_b_id_ex_int[9] , \dp/op_b_id_ex_int[8] ,
         \dp/op_b_id_ex_int[7] , \dp/op_b_id_ex_int[6] ,
         \dp/op_b_id_ex_int[5] , \dp/op_b_id_ex_int[4] ,
         \dp/op_b_id_ex_int[3] , \dp/op_b_id_ex_int[2] ,
         \dp/op_b_id_ex_int[1] , \dp/op_b_id_ex_int[0] , \dp/imm_id_int[15] ,
         \dp/imm_id_int[14] , \dp/imm_id_int[13] , \dp/imm_id_int[12] ,
         \dp/imm_id_int[11] , \dp/imm_id_int[10] , \dp/imm_id_int[9] ,
         \dp/imm_id_int[8] , \dp/imm_id_int[7] , \dp/imm_id_int[6] ,
         \dp/imm_id_int[5] , \dp/imm_id_int[4] , \dp/imm_id_int[3] ,
         \dp/imm_id_int[2] , \dp/imm_id_int[1] , \dp/imm_id_int[0] ,
         \dp/alu_out_low_mem_wb_int[0] , \dp/alu_out_low_mem_wb_int[1] ,
         \dp/alu_out_low_mem_wb_int[2] , \dp/alu_out_low_mem_wb_int[3] ,
         \dp/alu_out_low_mem_wb_int[4] , \dp/alu_out_low_mem_wb_int[5] ,
         \dp/alu_out_low_mem_wb_int[6] , \dp/alu_out_low_mem_wb_int[7] ,
         \dp/alu_out_low_mem_wb_int[8] , \dp/alu_out_low_mem_wb_int[9] ,
         \dp/alu_out_low_mem_wb_int[10] , \dp/alu_out_low_mem_wb_int[11] ,
         \dp/alu_out_low_mem_wb_int[12] , \dp/alu_out_low_mem_wb_int[13] ,
         \dp/alu_out_low_mem_wb_int[14] , \dp/alu_out_low_mem_wb_int[15] ,
         \dp/alu_out_low_mem_wb_int[16] , \dp/alu_out_low_mem_wb_int[17] ,
         \dp/alu_out_low_mem_wb_int[18] , \dp/alu_out_low_mem_wb_int[19] ,
         \dp/alu_out_low_mem_wb_int[20] , \dp/alu_out_low_mem_wb_int[21] ,
         \dp/alu_out_low_mem_wb_int[22] , \dp/alu_out_low_mem_wb_int[23] ,
         \dp/alu_out_low_mem_wb_int[24] , \dp/alu_out_low_mem_wb_int[25] ,
         \dp/alu_out_low_mem_wb_int[26] , \dp/alu_out_low_mem_wb_int[27] ,
         \dp/alu_out_low_mem_wb_int[28] , \dp/alu_out_low_mem_wb_int[29] ,
         \dp/alu_out_low_mem_wb_int[30] , \dp/alu_out_low_mem_wb_int[31] ,
         \dp/npc_id_exe_int[2] , \dp/npc_id_exe_int[3] ,
         \dp/npc_id_exe_int[4] , \dp/npc_id_exe_int[5] ,
         \dp/npc_id_exe_int[6] , \dp/npc_id_exe_int[7] ,
         \dp/npc_id_exe_int[8] , \dp/npc_id_exe_int[10] ,
         \dp/npc_id_exe_int[12] , \dp/npc_id_exe_int[14] ,
         \dp/npc_id_exe_int[16] , \dp/npc_id_exe_int[17] ,
         \dp/npc_id_exe_int[18] , \dp/npc_id_exe_int[20] ,
         \dp/npc_id_exe_int[21] , \dp/npc_id_exe_int[22] ,
         \dp/npc_id_exe_int[23] , \dp/npc_id_exe_int[24] ,
         \dp/npc_id_exe_int[25] , \dp/npc_id_exe_int[26] ,
         \dp/npc_id_exe_int[28] , \dp/npc_id_exe_int[31] ,
         \dp/pc_plus4_out_if_int[28] , \dp/pc_plus4_out_if_int[27] ,
         \dp/pc_plus4_out_if_int[26] , \dp/pc_plus4_out_if_int[25] ,
         \dp/pc_plus4_out_if_int[24] , \dp/pc_plus4_out_if_int[23] ,
         \dp/pc_plus4_out_if_int[22] , \dp/pc_plus4_out_if_int[21] ,
         \dp/pc_plus4_out_if_int[20] , \dp/pc_plus4_out_if_int[19] ,
         \dp/pc_plus4_out_if_int[18] , \dp/pc_plus4_out_if_int[17] ,
         \dp/pc_plus4_out_if_int[16] , \dp/pc_plus4_out_if_int[15] ,
         \dp/pc_plus4_out_if_int[14] , \dp/pc_plus4_out_if_int[13] ,
         \dp/pc_plus4_out_if_int[12] , \dp/pc_plus4_out_if_int[11] ,
         \dp/pc_plus4_out_if_int[10] , \dp/pc_plus4_out_if_int[9] ,
         \dp/pc_plus4_out_if_int[8] , \dp/pc_plus4_out_if_int[7] ,
         \dp/pc_plus4_out_if_int[6] , \dp/pc_plus4_out_if_int[5] ,
         \dp/pc_plus4_out_if_int[4] , \dp/pc_plus4_out_if_int[3] ,
         \dp/pc_plus4_out_if_int[2] , \dp/pc_plus4_out_if_int[1] ,
         \mc/currstate[0] , \mc/currstate[1] , \dp/ifs/pc_btb[29] ,
         \dp/ifs/pc_btb[28] , \dp/ifs/pc_btb[27] , \dp/ifs/pc_btb[26] ,
         \dp/ifs/pc_btb[25] , \dp/ifs/pc_btb[24] , \dp/ifs/pc_btb[23] ,
         \dp/ifs/pc_btb[22] , \dp/ifs/pc_btb[21] , \dp/ifs/pc_btb[20] ,
         \dp/ifs/pc_btb[19] , \dp/ifs/pc_btb[18] , \dp/ifs/pc_btb[17] ,
         \dp/ifs/pc_btb[16] , \dp/ifs/pc_btb[15] , \dp/ifs/pc_btb[14] ,
         \dp/ifs/pc_btb[13] , \dp/ifs/pc_btb[12] , \dp/ifs/pc_btb[11] ,
         \dp/ifs/pc_btb[10] , \dp/ifs/pc_btb[9] , \dp/ifs/pc_btb[8] ,
         \dp/ifs/pc_btb[7] , \dp/ifs/pc_btb[6] , \dp/ifs/pc_btb[5] ,
         \dp/ifs/pc_btb[4] , \dp/ifs/pc_btb[3] , \dp/ifs/pc_btb[2] ,
         \dp/ifs/pc_btb[1] , \dp/ifs/pc_btb[0] , \dp/ids/rp2[0] ,
         \dp/ids/rp2[1] , \dp/ids/rp2[2] , \dp/ids/rp2[3] , \dp/ids/rp2[4] ,
         \dp/ids/rp2[5] , \dp/ids/rp2[6] , \dp/ids/rp2[7] , \dp/ids/rp2[8] ,
         \dp/ids/rp2[9] , \dp/ids/rp2[10] , \dp/ids/rp2[11] , \dp/ids/rp2[12] ,
         \dp/ids/rp2[13] , \dp/ids/rp2[14] , \dp/ids/rp2[15] ,
         \dp/ids/rp2[16] , \dp/ids/rp2[17] , \dp/ids/rp2[18] ,
         \dp/ids/rp2[19] , \dp/ids/rp2[20] , \dp/ids/rp2[21] ,
         \dp/ids/rp2[22] , \dp/ids/rp2[23] , \dp/ids/rp2[24] ,
         \dp/ids/rp2[25] , \dp/ids/rp2[26] , \dp/ids/rp2[27] ,
         \dp/ids/rp2[28] , \dp/ids/rp2[29] , \dp/ids/rp2[30] ,
         \dp/ids/rp2[31] , \dp/ids/rp1[31] , \dp/ids/rp1[30] ,
         \dp/ids/rp1[29] , \dp/ids/rp1[28] , \dp/ids/rp1[27] ,
         \dp/ids/rp1[26] , \dp/ids/rp1[25] , \dp/ids/rp1[24] ,
         \dp/ids/rp1[23] , \dp/ids/rp1[22] , \dp/ids/rp1[21] ,
         \dp/ids/rp1[20] , \dp/ids/rp1[19] , \dp/ids/rp1[18] ,
         \dp/ids/rp1[17] , \dp/ids/rp1[16] , \dp/ids/rp1[15] ,
         \dp/ids/rp1[14] , \dp/ids/rp1[13] , \dp/ids/rp1[12] ,
         \dp/ids/rp1[11] , \dp/ids/rp1[10] , \dp/ids/rp1[9] , \dp/ids/rp1[8] ,
         \dp/ids/rp1[7] , \dp/ids/rp1[6] , \dp/ids/rp1[5] , \dp/ids/rp1[4] ,
         \dp/ids/rp1[3] , \dp/ids/rp1[2] , \dp/ids/rp1[1] , \dp/ids/rp1[0] ,
         \dp/exs/a_shift_int[31] , \dp/exs/a_shift_int[30] ,
         \dp/exs/a_shift_int[29] , \dp/exs/a_shift_int[28] ,
         \dp/exs/a_shift_int[27] , \dp/exs/a_shift_int[26] ,
         \dp/exs/a_shift_int[25] , \dp/exs/a_shift_int[24] ,
         \dp/exs/a_shift_int[23] , \dp/exs/a_shift_int[22] ,
         \dp/exs/a_shift_int[21] , \dp/exs/a_shift_int[20] ,
         \dp/exs/a_shift_int[19] , \dp/exs/a_shift_int[18] ,
         \dp/exs/a_shift_int[17] , \dp/exs/a_shift_int[16] ,
         \dp/exs/a_shift_int[15] , \dp/exs/a_shift_int[14] ,
         \dp/exs/a_shift_int[13] , \dp/exs/a_shift_int[12] ,
         \dp/exs/a_shift_int[11] , \dp/exs/a_shift_int[10] ,
         \dp/exs/a_shift_int[9] , \dp/exs/a_shift_int[8] ,
         \dp/exs/a_shift_int[7] , \dp/exs/a_shift_int[6] ,
         \dp/exs/a_shift_int[5] , \dp/exs/a_shift_int[4] ,
         \dp/exs/a_shift_int[3] , \dp/exs/a_shift_int[2] ,
         \dp/exs/a_shift_int[1] , \dp/exs/a_shift_int[0] ,
         \dp/id_exe_regs/b_mult_reg/q[17] , \dp/id_exe_regs/b_mult_reg/q[18] ,
         \dp/id_exe_regs/b_mult_reg/q[19] , \dp/id_exe_regs/b_mult_reg/q[20] ,
         \dp/id_exe_regs/b_mult_reg/q[21] , \dp/id_exe_regs/b_mult_reg/q[22] ,
         \dp/id_exe_regs/b_mult_reg/q[23] , \dp/id_exe_regs/b_mult_reg/q[24] ,
         \dp/id_exe_regs/b_mult_reg/q[25] , \dp/id_exe_regs/b_mult_reg/q[26] ,
         \dp/id_exe_regs/b_mult_reg/q[27] , \dp/id_exe_regs/b_mult_reg/q[28] ,
         \dp/id_exe_regs/b_mult_reg/q[29] , \dp/id_exe_regs/b_mult_reg/q[30] ,
         \dp/exs/alu_unit/shifter_out[31] , \dp/exs/alu_unit/shifter_out[30] ,
         \dp/exs/alu_unit/shifter_out[29] , \dp/exs/alu_unit/shifter_out[28] ,
         \dp/exs/alu_unit/shifter_out[27] , \dp/exs/alu_unit/shifter_out[26] ,
         \dp/exs/alu_unit/shifter_out[25] , \dp/exs/alu_unit/shifter_out[24] ,
         \dp/exs/alu_unit/shifter_out[23] , \dp/exs/alu_unit/shifter_out[22] ,
         \dp/exs/alu_unit/shifter_out[21] , \dp/exs/alu_unit/shifter_out[20] ,
         \dp/exs/alu_unit/shifter_out[19] , \dp/exs/alu_unit/shifter_out[18] ,
         \dp/exs/alu_unit/shifter_out[17] , \dp/exs/alu_unit/shifter_out[16] ,
         \dp/exs/alu_unit/shifter_out[15] , \dp/exs/alu_unit/shifter_out[14] ,
         \dp/exs/alu_unit/shifter_out[13] , \dp/exs/alu_unit/shifter_out[12] ,
         \dp/exs/alu_unit/shifter_out[11] , \dp/exs/alu_unit/shifter_out[10] ,
         \dp/exs/alu_unit/shifter_out[9] , \dp/exs/alu_unit/shifter_out[8] ,
         \dp/exs/alu_unit/shifter_out[7] , \dp/exs/alu_unit/shifter_out[6] ,
         \dp/exs/alu_unit/shifter_out[5] , \dp/exs/alu_unit/shifter_out[4] ,
         \dp/exs/alu_unit/shifter_out[3] , \dp/exs/alu_unit/shifter_out[2] ,
         \dp/exs/alu_unit/shifter_out[1] , \dp/exs/alu_unit/shifter_out[0] ,
         \dp/exs/alu_unit/mult/neg_ax2_shiftn[12] ,
         \dp/exs/alu_unit/mult/neg_ax2_shiftn[11] ,
         \dp/exs/alu_unit/mult/neg_ax2_shiftn[10] ,
         \dp/exs/alu_unit/mult/neg_ax2_shiftn[9] ,
         \dp/exs/alu_unit/mult/neg_ax2_shiftn[8] ,
         \dp/exs/alu_unit/mult/neg_ax2_shiftn[7] ,
         \dp/exs/alu_unit/mult/neg_ax2_shiftn[6] ,
         \dp/exs/alu_unit/mult/neg_ax2_shiftn[5] ,
         \dp/exs/alu_unit/mult/neg_ax2_shiftn[4] ,
         \dp/exs/alu_unit/mult/ax2_shiftn[12] ,
         \dp/exs/alu_unit/mult/ax2_shiftn[11] ,
         \dp/exs/alu_unit/mult/ax2_shiftn[10] ,
         \dp/exs/alu_unit/mult/ax2_shiftn[9] ,
         \dp/exs/alu_unit/mult/ax2_shiftn[8] ,
         \dp/exs/alu_unit/mult/ax2_shiftn[7] ,
         \dp/exs/alu_unit/mult/ax2_shiftn[6] ,
         \dp/exs/alu_unit/mult/ax2_shiftn[5] ,
         \dp/exs/alu_unit/mult/ax2_shiftn[4] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[63] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[62] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[61] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[60] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[59] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[58] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[57] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[56] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[55] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[54] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[53] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[52] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[51] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[50] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[49] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[48] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[47] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[46] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[45] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[44] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[43] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[42] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[41] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[40] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[39] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[38] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[37] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[36] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[35] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[34] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[33] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[32] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[31] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[30] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[29] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[28] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[27] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[26] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[25] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[24] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[23] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[22] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[21] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[20] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[19] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[18] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[17] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[16] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[15] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[14] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[13] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[12] ,
         \dp/exs/alu_unit/mult/neg_a_shiftn[2] ,
         \dp/exs/alu_unit/mult/a_shiftn[63] ,
         \dp/exs/alu_unit/mult/a_shiftn[62] ,
         \dp/exs/alu_unit/mult/a_shiftn[61] ,
         \dp/exs/alu_unit/mult/a_shiftn[60] ,
         \dp/exs/alu_unit/mult/a_shiftn[59] ,
         \dp/exs/alu_unit/mult/a_shiftn[58] ,
         \dp/exs/alu_unit/mult/a_shiftn[57] ,
         \dp/exs/alu_unit/mult/a_shiftn[56] ,
         \dp/exs/alu_unit/mult/a_shiftn[55] ,
         \dp/exs/alu_unit/mult/a_shiftn[54] ,
         \dp/exs/alu_unit/mult/a_shiftn[53] ,
         \dp/exs/alu_unit/mult/a_shiftn[52] ,
         \dp/exs/alu_unit/mult/a_shiftn[51] ,
         \dp/exs/alu_unit/mult/a_shiftn[50] ,
         \dp/exs/alu_unit/mult/a_shiftn[49] ,
         \dp/exs/alu_unit/mult/a_shiftn[48] ,
         \dp/exs/alu_unit/mult/a_shiftn[47] ,
         \dp/exs/alu_unit/mult/a_shiftn[46] ,
         \dp/exs/alu_unit/mult/a_shiftn[45] ,
         \dp/exs/alu_unit/mult/a_shiftn[44] ,
         \dp/exs/alu_unit/mult/a_shiftn[43] ,
         \dp/exs/alu_unit/mult/a_shiftn[42] ,
         \dp/exs/alu_unit/mult/a_shiftn[41] ,
         \dp/exs/alu_unit/mult/a_shiftn[40] ,
         \dp/exs/alu_unit/mult/a_shiftn[39] ,
         \dp/exs/alu_unit/mult/a_shiftn[38] ,
         \dp/exs/alu_unit/mult/a_shiftn[37] ,
         \dp/exs/alu_unit/mult/a_shiftn[36] ,
         \dp/exs/alu_unit/mult/a_shiftn[35] ,
         \dp/exs/alu_unit/mult/a_shiftn[34] ,
         \dp/exs/alu_unit/mult/a_shiftn[33] ,
         \dp/exs/alu_unit/mult/a_shiftn[32] ,
         \dp/exs/alu_unit/mult/a_shiftn[31] ,
         \dp/exs/alu_unit/mult/a_shiftn[30] ,
         \dp/exs/alu_unit/mult/a_shiftn[29] ,
         \dp/exs/alu_unit/mult/a_shiftn[28] ,
         \dp/exs/alu_unit/mult/a_shiftn[27] ,
         \dp/exs/alu_unit/mult/a_shiftn[26] ,
         \dp/exs/alu_unit/mult/a_shiftn[25] ,
         \dp/exs/alu_unit/mult/a_shiftn[24] ,
         \dp/exs/alu_unit/mult/a_shiftn[23] ,
         \dp/exs/alu_unit/mult/a_shiftn[22] ,
         \dp/exs/alu_unit/mult/a_shiftn[21] ,
         \dp/exs/alu_unit/mult/a_shiftn[20] ,
         \dp/exs/alu_unit/mult/a_shiftn[19] ,
         \dp/exs/alu_unit/mult/a_shiftn[18] ,
         \dp/exs/alu_unit/mult/a_shiftn[17] ,
         \dp/exs/alu_unit/mult/a_shiftn[16] ,
         \dp/exs/alu_unit/mult/a_shiftn[15] ,
         \dp/exs/alu_unit/mult/a_shiftn[14] ,
         \dp/exs/alu_unit/mult/a_shiftn[13] ,
         \dp/exs/alu_unit/mult/a_shiftn[12] ,
         \dp/exs/alu_unit/mult/a_shiftn[2] , n92, n95, n99, n103, n110, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n288, n289, n290, n291, n292, n293, n294, n295, n299, n300,
         n301, n302, n303, n304, n305, n306, n307, n308, n309, n310, n311,
         n312, n313, n314, n315, n316, n317, n318, n319, n320, n321, n322,
         n323, n324, n325, n326, n327, n328, n329, n330, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n463, n465, n466, n467, n471, n472,
         n473, n474, n478, n479, n480, n490, n491, n492, n493, n494, n593,
         n594, n595, n613, n614, n615, n616, n617, n618, n619, n620, n621,
         n622, n623, n624, n625, n626, n627, n628, n629, n630, n631, n632,
         n633, n634, n635, n636, n637, n638, n639, n640, n641, n642, n643,
         n644, n681, n1143, n1144, n1444, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1493, n1594, n1597, n1598, n1599,
         n1600, n1603, n1604, n1605, n1606, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2725, n2726, n2727, n2728, n2729,
         n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909,
         n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919,
         n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929,
         n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939,
         n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949,
         n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959,
         n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989,
         n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999,
         n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, \ctrl_u/n560 ,
         \ctrl_u/n559 , \ctrl_u/n558 , \ctrl_u/n557 , \ctrl_u/n556 ,
         \ctrl_u/n555 , \ctrl_u/n554 , \ctrl_u/n553 , \ctrl_u/n552 ,
         \ctrl_u/n551 , \ctrl_u/n550 , \ctrl_u/n549 , \ctrl_u/n548 ,
         \ctrl_u/n547 , \ctrl_u/n546 , \ctrl_u/n545 , \ctrl_u/n544 ,
         \ctrl_u/n543 , \ctrl_u/n542 , \ctrl_u/n541 , \ctrl_u/n540 ,
         \ctrl_u/n539 , \ctrl_u/n538 , \ctrl_u/n537 , \ctrl_u/n536 ,
         \ctrl_u/n535 , \ctrl_u/n534 , \ctrl_u/n533 , \ctrl_u/n532 ,
         \ctrl_u/n531 , \ctrl_u/n530 , \ctrl_u/n528 , \ctrl_u/n527 ,
         \ctrl_u/n526 , \ctrl_u/n524 , \ctrl_u/n523 , \ctrl_u/n522 ,
         \ctrl_u/n521 , \ctrl_u/n520 , \ctrl_u/n519 , \ctrl_u/n518 ,
         \ctrl_u/n517 , \ctrl_u/n514 , \ctrl_u/n513 , \ctrl_u/n512 ,
         \ctrl_u/n511 , \ctrl_u/n510 , \ctrl_u/n509 , \ctrl_u/n508 ,
         \ctrl_u/n507 , \ctrl_u/n506 , \ctrl_u/n505 , \ctrl_u/n504 ,
         \ctrl_u/n503 , \ctrl_u/n502 , \ctrl_u/n501 , \ctrl_u/n486 ,
         \ctrl_u/n484 , \ctrl_u/n483 , \ctrl_u/n481 , \ctrl_u/n480 ,
         \ctrl_u/n479 , \ctrl_u/n478 , \ctrl_u/n477 , \ctrl_u/n476 ,
         \ctrl_u/n475 , \ctrl_u/n474 , \ctrl_u/n473 , \ctrl_u/n472 ,
         \ctrl_u/n471 , \ctrl_u/n470 , \ctrl_u/n469 , \ctrl_u/n468 ,
         \ctrl_u/n467 , \ctrl_u/n465 , \ctrl_u/n461 , \ctrl_u/n460 ,
         \ctrl_u/n459 , \ctrl_u/n458 , \ctrl_u/n457 , \ctrl_u/n456 ,
         \ctrl_u/n455 , \ctrl_u/n454 , \ctrl_u/n453 , \ctrl_u/n452 ,
         \ctrl_u/n451 , \ctrl_u/n450 , \ctrl_u/n449 , \ctrl_u/n448 ,
         \ctrl_u/n447 , \ctrl_u/n446 , \ctrl_u/n445 , \ctrl_u/n444 ,
         \ctrl_u/n443 , \ctrl_u/n442 , \ctrl_u/n441 , \ctrl_u/n440 ,
         \ctrl_u/n439 , \ctrl_u/n438 , \ctrl_u/n437 , \ctrl_u/n436 ,
         \ctrl_u/n435 , \ctrl_u/n434 , \ctrl_u/n433 , \ctrl_u/n432 ,
         \ctrl_u/n430 , \ctrl_u/n429 , \ctrl_u/n428 , \ctrl_u/n427 ,
         \ctrl_u/n426 , \ctrl_u/n425 , \ctrl_u/n423 , \ctrl_u/n422 ,
         \ctrl_u/n421 , \ctrl_u/n420 , \ctrl_u/n412 , \ctrl_u/n406 ,
         \ctrl_u/n402 , \ctrl_u/n386 , \ctrl_u/n384 , \ctrl_u/n335 ,
         \ctrl_u/n305 , \ctrl_u/n303 , \ctrl_u/n301 , \ctrl_u/n245 ,
         \ctrl_u/n193 , \ctrl_u/n181 , \ctrl_u/n179 , \ctrl_u/n170 ,
         \ctrl_u/n169 , \ctrl_u/n167 , \ctrl_u/n166 , \ctrl_u/n95 ,
         \ctrl_u/n94 , \ctrl_u/n83 , \ctrl_u/n74 , \ctrl_u/n73 , \ctrl_u/n72 ,
         \ctrl_u/n70 , \ctrl_u/n69 , \ctrl_u/n68 , \ctrl_u/n67 , \ctrl_u/n66 ,
         \ctrl_u/n65 , \ctrl_u/n64 , \ctrl_u/n63 , \ctrl_u/n62 , \ctrl_u/n61 ,
         \ctrl_u/n59 , \ctrl_u/n27 , \ctrl_u/n25 , \ctrl_u/n23 , \ctrl_u/n21 ,
         \ctrl_u/n15 , \ctrl_u/n13 , \ctrl_u/n11 , \ctrl_u/n9 , \ctrl_u/N1805 ,
         \ctrl_u/mem_stall , \ctrl_u/exe_stall , \ctrl_u/if_stall ,
         \ctrl_u/next_mem[10] , \ctrl_u/next_mem[8] , \ctrl_u/next_mem[7] ,
         \ctrl_u/next_mem[6] , \ctrl_u/next_mem[4] , \ctrl_u/next_mem[3] ,
         \ctrl_u/next_mem[2] , \ctrl_u/curr_mul_end_wb ,
         \ctrl_u/curr_mul_end_mem , \ctrl_u/curr_ms , \ctrl_u/curr_wb[3] ,
         \ctrl_u/curr_mem[0] , \ctrl_u/curr_mem[1] , \ctrl_u/curr_mem[2] ,
         \ctrl_u/curr_mem[3] , \ctrl_u/curr_mem[4] , \ctrl_u/curr_mem[5] ,
         \ctrl_u/curr_mem[6] , \ctrl_u/curr_mem_11 , \ctrl_u/curr_mem_12 ,
         \ctrl_u/next_exe[41] , \ctrl_u/next_exe[40] , \ctrl_u/next_exe[39] ,
         \ctrl_u/next_exe[38] , \ctrl_u/next_exe[36] , \ctrl_u/next_exe[33] ,
         \ctrl_u/next_exe[32] , \ctrl_u/next_exe[31] , \ctrl_u/next_exe[28] ,
         \ctrl_u/next_exe[27] , \ctrl_u/next_exe[21] , \ctrl_u/next_exe[20] ,
         \ctrl_u/next_exe[19] , \ctrl_u/next_exe[16] , \ctrl_u/next_exe[14] ,
         \ctrl_u/next_exe[13] , \ctrl_u/next_exe[12] , \ctrl_u/next_exe[11] ,
         \ctrl_u/next_exe[10] , \ctrl_u/next_exe[9] , \ctrl_u/next_exe[8] ,
         \ctrl_u/next_exe[7] , \ctrl_u/next_exe[5] , \ctrl_u/next_exe[1] ,
         \ctrl_u/next_exe[0] , \ctrl_u/curr_mul_in_prog , \ctrl_u/curr_pt_exe ,
         \ctrl_u/curr_ak_exe , \ctrl_u/curr_exe[0] , \ctrl_u/curr_exe[1] ,
         \ctrl_u/curr_exe[2] , \ctrl_u/curr_exe[3] , \ctrl_u/curr_exe[4] ,
         \ctrl_u/curr_exe[5] , \ctrl_u/curr_exe[6] , \ctrl_u/curr_exe[7] ,
         \ctrl_u/curr_exe[8] , \ctrl_u/curr_exe[9] , \ctrl_u/curr_exe[10] ,
         \ctrl_u/curr_exe[11] , \ctrl_u/curr_exe[12] , \ctrl_u/curr_exe[13] ,
         \ctrl_u/curr_exe[14] , \ctrl_u/curr_exe[15] , \ctrl_u/curr_exe[16] ,
         \ctrl_u/curr_exe[17] , \ctrl_u/curr_exe[18] , \ctrl_u/curr_exe[19] ,
         \ctrl_u/curr_exe[20] , \ctrl_u/curr_exe_39 , \ctrl_u/curr_exe_40 ,
         \ctrl_u/curr_exe_41 , \ctrl_u/curr_pt_id , \ctrl_u/curr_ak_id ,
         \ctrl_u/curr_id[0] , \ctrl_u/curr_id[1] , \ctrl_u/curr_id[2] ,
         \ctrl_u/curr_id[3] , \ctrl_u/curr_id[4] , \ctrl_u/curr_id[5] ,
         \ctrl_u/curr_id[6] , \ctrl_u/curr_id[7] , \ctrl_u/curr_id[8] ,
         \ctrl_u/curr_id[9] , \ctrl_u/curr_id[10] , \ctrl_u/curr_id[11] ,
         \ctrl_u/curr_id[12] , \ctrl_u/curr_id[13] , \ctrl_u/curr_id[14] ,
         \ctrl_u/curr_id[16] , \ctrl_u/curr_id[17] , \ctrl_u/curr_id[18] ,
         \ctrl_u/curr_id[19] , \ctrl_u/curr_id[20] , \ctrl_u/curr_id[21] ,
         \ctrl_u/curr_id[22] , \ctrl_u/curr_id[25] , \ctrl_u/curr_id[26] ,
         \ctrl_u/curr_id[27] , \ctrl_u/curr_id[28] , \ctrl_u/curr_id[29] ,
         \ctrl_u/curr_id[31] , \ctrl_u/curr_id[32] , \ctrl_u/curr_id[33] ,
         \ctrl_u/curr_id[34] , \ctrl_u/curr_id[35] , \ctrl_u/curr_id[36] ,
         \ctrl_u/curr_id[38] , \ctrl_u/curr_id[39] , \ctrl_u/curr_id[40] ,
         \ctrl_u/curr_id[41] , \ctrl_u/op_type_exe[1] , \intadd_2/A[8] ,
         \intadd_2/A[6] , \intadd_2/A[4] , \intadd_2/A[2] , \intadd_2/A[0] ,
         \intadd_2/B[20] , \intadd_2/B[14] , \intadd_2/SUM[27] ,
         \intadd_2/SUM[26] , \intadd_2/SUM[25] , \intadd_2/SUM[24] ,
         \intadd_2/SUM[23] , \intadd_2/SUM[22] , \intadd_2/SUM[21] ,
         \intadd_2/SUM[20] , \intadd_2/SUM[19] , \intadd_2/SUM[18] ,
         \intadd_2/SUM[17] , \intadd_2/SUM[16] , \intadd_2/SUM[15] ,
         \intadd_2/SUM[14] , \intadd_2/SUM[13] , \intadd_2/SUM[12] ,
         \intadd_2/SUM[11] , \intadd_2/SUM[10] , \intadd_2/SUM[9] ,
         \intadd_2/SUM[8] , \intadd_2/SUM[7] , \intadd_2/SUM[6] ,
         \intadd_2/SUM[5] , \intadd_2/SUM[4] , \intadd_2/SUM[3] ,
         \intadd_2/SUM[2] , \intadd_2/SUM[1] , \intadd_2/SUM[0] ,
         \intadd_2/n23 , \intadd_2/n22 , \intadd_2/n21 , \intadd_2/n20 ,
         \intadd_2/n19 , \intadd_2/n18 , \intadd_2/n17 , \intadd_2/n13 ,
         \intadd_2/n12 , \intadd_2/n11 , \intadd_2/n6 , \intadd_2/n5 ,
         \intadd_2/n4 , \intadd_2/n3 , \intadd_2/n2 , \intadd_1/A[29] ,
         \intadd_1/A[28] , \intadd_1/A[27] , \intadd_1/A[26] ,
         \intadd_1/A[25] , \intadd_1/A[24] , \intadd_1/A[23] ,
         \intadd_1/A[21] , \intadd_1/A[19] , \intadd_1/A[18] ,
         \intadd_1/A[17] , \intadd_1/A[16] , \intadd_1/A[15] ,
         \intadd_1/A[14] , \intadd_1/A[13] , \intadd_1/A[12] ,
         \intadd_1/A[11] , \intadd_1/A[9] , \intadd_1/A[8] , \intadd_1/A[7] ,
         \intadd_1/A[6] , \intadd_1/A[5] , \intadd_1/A[3] , \intadd_1/A[2] ,
         \intadd_1/A[1] , \intadd_1/A[0] , \intadd_1/B[29] , \intadd_1/B[28] ,
         \intadd_1/B[27] , \intadd_1/B[26] , \intadd_1/B[25] ,
         \intadd_1/B[24] , \intadd_1/B[23] , \intadd_1/B[22] ,
         \intadd_1/B[21] , \intadd_1/B[20] , \intadd_1/B[19] ,
         \intadd_1/B[18] , \intadd_1/B[17] , \intadd_1/B[16] ,
         \intadd_1/B[15] , \intadd_1/B[14] , \intadd_1/B[13] ,
         \intadd_1/B[12] , \intadd_1/B[11] , \intadd_1/B[10] , \intadd_1/B[9] ,
         \intadd_1/B[8] , \intadd_1/B[7] , \intadd_1/B[6] , \intadd_1/B[5] ,
         \intadd_1/B[4] , \intadd_1/B[3] , \intadd_1/B[2] , \intadd_1/B[1] ,
         \intadd_1/B[0] , \intadd_1/CI , \intadd_1/SUM[29] ,
         \intadd_1/SUM[28] , \intadd_1/SUM[27] , \intadd_1/SUM[26] ,
         \intadd_1/SUM[25] , \intadd_1/SUM[24] , \intadd_1/SUM[23] ,
         \intadd_1/SUM[22] , \intadd_1/SUM[21] , \intadd_1/SUM[20] ,
         \intadd_1/SUM[19] , \intadd_1/SUM[18] , \intadd_1/SUM[17] ,
         \intadd_1/SUM[16] , \intadd_1/SUM[15] , \intadd_1/SUM[14] ,
         \intadd_1/SUM[13] , \intadd_1/SUM[12] , \intadd_1/SUM[11] ,
         \intadd_1/SUM[10] , \intadd_1/SUM[9] , \intadd_1/SUM[8] ,
         \intadd_1/SUM[7] , \intadd_1/SUM[6] , \intadd_1/SUM[5] ,
         \intadd_1/SUM[3] , \intadd_1/SUM[2] , \intadd_1/SUM[1] ,
         \intadd_1/SUM[0] , \intadd_1/n199 , \intadd_1/n198 , \intadd_1/n196 ,
         \intadd_1/n193 , \intadd_1/n192 , \intadd_1/n191 , \intadd_1/n190 ,
         \intadd_1/n188 , \intadd_1/n186 , \intadd_1/n185 , \intadd_1/n183 ,
         \intadd_1/n182 , \intadd_1/n181 , \intadd_1/n179 , \intadd_1/n177 ,
         \intadd_1/n173 , \intadd_1/n172 , \intadd_1/n171 , \intadd_1/n169 ,
         \intadd_1/n168 , \intadd_1/n167 , \intadd_1/n166 , \intadd_1/n165 ,
         \intadd_1/n164 , \intadd_1/n163 , \intadd_1/n162 , \intadd_1/n161 ,
         \intadd_1/n160 , \intadd_1/n159 , \intadd_1/n158 , \intadd_1/n154 ,
         \intadd_1/n153 , \intadd_1/n152 , \intadd_1/n151 , \intadd_1/n150 ,
         \intadd_1/n149 , \intadd_1/n148 , \intadd_1/n147 , \intadd_1/n146 ,
         \intadd_1/n145 , \intadd_1/n144 , \intadd_1/n143 , \intadd_1/n142 ,
         \intadd_1/n141 , \intadd_1/n140 , \intadd_1/n139 , \intadd_1/n138 ,
         \intadd_1/n137 , \intadd_1/n136 , \intadd_1/n135 , \intadd_1/n134 ,
         \intadd_1/n132 , \intadd_1/n131 , \intadd_1/n130 , \intadd_1/n128 ,
         \intadd_1/n127 , \intadd_1/n123 , \intadd_1/n122 , \intadd_1/n121 ,
         \intadd_1/n120 , \intadd_1/n119 , \intadd_1/n118 , \intadd_1/n117 ,
         \intadd_1/n115 , \intadd_1/n114 , \intadd_1/n113 , \intadd_1/n111 ,
         \intadd_1/n110 , \intadd_1/n109 , \intadd_1/n108 , \intadd_1/n107 ,
         \intadd_1/n104 , \intadd_1/n103 , \intadd_1/n102 , \intadd_1/n101 ,
         \intadd_1/n99 , \intadd_1/n98 , \intadd_1/n97 , \intadd_1/n96 ,
         \intadd_1/n95 , \intadd_1/n94 , \intadd_1/n93 , \intadd_1/n92 ,
         \intadd_1/n91 , \intadd_1/n90 , \intadd_1/n89 , \intadd_1/n88 ,
         \intadd_1/n87 , \intadd_1/n86 , \intadd_1/n85 , \intadd_1/n84 ,
         \intadd_1/n83 , \intadd_1/n82 , \intadd_1/n81 , \intadd_1/n80 ,
         \intadd_1/n78 , \intadd_1/n77 , \intadd_1/n75 , \intadd_1/n74 ,
         \intadd_1/n73 , \intadd_1/n72 , \intadd_1/n71 , \intadd_1/n70 ,
         \intadd_1/n69 , \intadd_1/n68 , \intadd_1/n65 , \intadd_1/n64 ,
         \intadd_1/n63 , \intadd_1/n62 , \intadd_1/n61 , \intadd_1/n60 ,
         \intadd_1/n59 , \intadd_1/n57 , \intadd_1/n56 , \intadd_1/n55 ,
         \intadd_1/n54 , \intadd_1/n53 , \intadd_1/n52 , \intadd_1/n51 ,
         \intadd_1/n50 , \intadd_1/n49 , \intadd_1/n48 , \intadd_1/n47 ,
         \intadd_1/n46 , \intadd_1/n45 , \intadd_1/n43 , \intadd_1/n41 ,
         \intadd_1/n40 , \intadd_1/n39 , \intadd_1/n38 , \intadd_1/n37 ,
         \intadd_1/n36 , \intadd_1/n33 , \intadd_1/n30 , \intadd_1/n28 ,
         \intadd_1/n26 , \intadd_1/n25 , \intadd_1/n24 , \intadd_1/n23 ,
         \intadd_1/n20 , \intadd_1/n19 , \intadd_1/n18 , \intadd_1/n17 ,
         \intadd_1/n15 , \intadd_1/n14 , \intadd_1/n13 , \intadd_1/n12 ,
         \intadd_1/n11 , \intadd_1/n8 , \intadd_1/n6 , \intadd_1/n4 ,
         \add_x_20/n28 , \add_x_20/n27 , \add_x_20/n26 , \add_x_20/n25 ,
         \add_x_20/n24 , \add_x_20/n23 , \add_x_20/n22 , \add_x_20/n21 ,
         \add_x_20/n20 , \add_x_20/n19 , \add_x_20/n18 , \add_x_20/n17 ,
         \add_x_20/n16 , \add_x_20/n15 , \add_x_20/n14 , \add_x_20/n13 ,
         \add_x_20/n12 , \add_x_20/n11 , \add_x_20/n10 , \add_x_20/n9 ,
         \add_x_20/n8 , \add_x_20/n7 , \add_x_20/n6 , \add_x_20/n5 ,
         \add_x_20/n4 , \add_x_20/n3 , \add_x_20/n2 , n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3970, n3974, n3975,
         n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983, n3984, n3985,
         n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993, n3994, n3995,
         n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003, n4004, n4005,
         n4007, n4008, n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016,
         n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026,
         n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036,
         n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046,
         n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056,
         n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106,
         n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116,
         n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126,
         n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136,
         n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146,
         n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156,
         n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166,
         n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176,
         n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186,
         n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196,
         n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206,
         n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216,
         n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226,
         n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236,
         n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246,
         n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256,
         n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266,
         n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276,
         n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286,
         n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296,
         n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306,
         n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316,
         n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326,
         n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336,
         n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346,
         n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356,
         n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366,
         n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376,
         n4377, n4378, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547,
         n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557,
         n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567,
         n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577,
         n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587,
         n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597,
         n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607,
         n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7264, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531;
  wire   [1:0] rp1_out_sel_id;
  wire   [1:0] rp2_out_sel_id;
  wire   [4:0] rs_id;
  wire   [4:0] rt_id;
  wire   [4:0] rd_idexe;
  wire   [3:0] shift_type_exe;
  wire   [3:0] log_type_exe;
  wire   [1:0] op_type_exe;
  wire   [3:0] it_exe;
  wire   [2:0] cond_sel_exe;
  wire   [2:0] alu_comp_sel;
  wire   [1:0] op_b_fw_sel_exe;
  wire   [4:0] rs_exe;
  wire   [4:0] rt_exe;
  wire   [4:0] rd_exemem;
  wire   [1:0] ld_type_mem;
  tri   dcache_update;
  tri   [1:0] dcache_update_type;
  tri   en_add_id;
  tri   en_mul_id;
  tri   en_shift_id;
  tri   en_a_neg_id;
  tri   shift_reg_id;
  tri   en_shift_reg_id;
  tri   en_rd_id;
  tri   en_npc_id;
  tri   en_imm_id;
  tri   en_b_id;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, 
        SYNOPSYS_UNCONNECTED__32, SYNOPSYS_UNCONNECTED__33, 
        SYNOPSYS_UNCONNECTED__34, SYNOPSYS_UNCONNECTED__35, 
        SYNOPSYS_UNCONNECTED__36, SYNOPSYS_UNCONNECTED__37, 
        SYNOPSYS_UNCONNECTED__38, SYNOPSYS_UNCONNECTED__39, 
        SYNOPSYS_UNCONNECTED__40, SYNOPSYS_UNCONNECTED__41, 
        SYNOPSYS_UNCONNECTED__42, SYNOPSYS_UNCONNECTED__43, 
        SYNOPSYS_UNCONNECTED__44, SYNOPSYS_UNCONNECTED__45, 
        SYNOPSYS_UNCONNECTED__46, SYNOPSYS_UNCONNECTED__47, 
        SYNOPSYS_UNCONNECTED__48, SYNOPSYS_UNCONNECTED__49, 
        SYNOPSYS_UNCONNECTED__50, SYNOPSYS_UNCONNECTED__51, 
        SYNOPSYS_UNCONNECTED__52, SYNOPSYS_UNCONNECTED__53, 
        SYNOPSYS_UNCONNECTED__54, SYNOPSYS_UNCONNECTED__55, 
        SYNOPSYS_UNCONNECTED__56, SYNOPSYS_UNCONNECTED__57, 
        SYNOPSYS_UNCONNECTED__58, SYNOPSYS_UNCONNECTED__59, 
        SYNOPSYS_UNCONNECTED__60, SYNOPSYS_UNCONNECTED__61, 
        SYNOPSYS_UNCONNECTED__62, SYNOPSYS_UNCONNECTED__63, 
        SYNOPSYS_UNCONNECTED__64, SYNOPSYS_UNCONNECTED__65, 
        SYNOPSYS_UNCONNECTED__66, SYNOPSYS_UNCONNECTED__67, 
        SYNOPSYS_UNCONNECTED__68, SYNOPSYS_UNCONNECTED__69, 
        SYNOPSYS_UNCONNECTED__70, SYNOPSYS_UNCONNECTED__71, 
        SYNOPSYS_UNCONNECTED__72, SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76, SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        SYNOPSYS_UNCONNECTED__128, SYNOPSYS_UNCONNECTED__129, 
        SYNOPSYS_UNCONNECTED__130, SYNOPSYS_UNCONNECTED__131;
  assign pc_out[29] = btb_cache_read_address[29];
  assign pc_out[28] = btb_cache_read_address[28];
  assign pc_out[27] = btb_cache_read_address[27];
  assign pc_out[26] = btb_cache_read_address[26];
  assign pc_out[25] = btb_cache_read_address[25];
  assign pc_out[24] = btb_cache_read_address[24];
  assign pc_out[23] = btb_cache_read_address[23];
  assign pc_out[22] = btb_cache_read_address[22];
  assign pc_out[21] = btb_cache_read_address[21];
  assign pc_out[20] = btb_cache_read_address[20];
  assign pc_out[19] = btb_cache_read_address[19];
  assign pc_out[18] = btb_cache_read_address[18];
  assign pc_out[17] = btb_cache_read_address[17];
  assign pc_out[16] = btb_cache_read_address[16];
  assign pc_out[15] = btb_cache_read_address[15];
  assign pc_out[14] = btb_cache_read_address[14];
  assign pc_out[13] = btb_cache_read_address[13];
  assign pc_out[12] = btb_cache_read_address[12];
  assign pc_out[11] = btb_cache_read_address[11];
  assign pc_out[10] = btb_cache_read_address[10];
  assign pc_out[9] = btb_cache_read_address[9];
  assign pc_out[8] = btb_cache_read_address[8];
  assign pc_out[7] = btb_cache_read_address[7];
  assign pc_out[6] = btb_cache_read_address[6];
  assign pc_out[5] = btb_cache_read_address[5];
  assign pc_out[4] = btb_cache_read_address[4];
  assign pc_out[3] = btb_cache_read_address[3];
  assign pc_out[2] = btb_cache_read_address[2];
  assign pc_out[1] = btb_cache_read_address[1];
  assign pc_out[0] = btb_cache_read_address[0];
  assign ram_to_cache_data[31] = ram_data_out[31];
  assign ram_to_cache_data[30] = ram_data_out[30];
  assign ram_to_cache_data[29] = ram_data_out[29];
  assign ram_to_cache_data[28] = ram_data_out[28];
  assign ram_to_cache_data[27] = ram_data_out[27];
  assign ram_to_cache_data[26] = ram_data_out[26];
  assign ram_to_cache_data[25] = ram_data_out[25];
  assign ram_to_cache_data[24] = ram_data_out[24];
  assign ram_to_cache_data[23] = ram_data_out[23];
  assign ram_to_cache_data[22] = ram_data_out[22];
  assign ram_to_cache_data[21] = ram_data_out[21];
  assign ram_to_cache_data[20] = ram_data_out[20];
  assign ram_to_cache_data[19] = ram_data_out[19];
  assign ram_to_cache_data[18] = ram_data_out[18];
  assign ram_to_cache_data[17] = ram_data_out[17];
  assign ram_to_cache_data[16] = ram_data_out[16];
  assign ram_to_cache_data[15] = ram_data_out[15];
  assign ram_to_cache_data[14] = ram_data_out[14];
  assign ram_to_cache_data[13] = ram_data_out[13];
  assign ram_to_cache_data[12] = ram_data_out[12];
  assign ram_to_cache_data[11] = ram_data_out[11];
  assign ram_to_cache_data[10] = ram_data_out[10];
  assign ram_to_cache_data[9] = ram_data_out[9];
  assign ram_to_cache_data[8] = ram_data_out[8];
  assign ram_to_cache_data[7] = ram_data_out[7];
  assign ram_to_cache_data[6] = ram_data_out[6];
  assign ram_to_cache_data[5] = ram_data_out[5];
  assign ram_to_cache_data[4] = ram_data_out[4];
  assign ram_to_cache_data[3] = ram_data_out[3];
  assign ram_to_cache_data[2] = ram_data_out[2];
  assign ram_to_cache_data[1] = ram_data_out[1];
  assign ram_to_cache_data[0] = ram_data_out[0];
  assign btb_addr_known_if = btb_cache_hit_read;
  assign rst_mem_wb_regs = rst;
  assign \dp/cache_in_mem_int[7]  = dcache_data_in[7];
  assign \dp/cache_in_mem_int[6]  = dcache_data_in[6];
  assign \dp/cache_in_mem_int[5]  = dcache_data_in[5];
  assign \dp/cache_in_mem_int[4]  = dcache_data_in[4];
  assign \dp/cache_in_mem_int[3]  = dcache_data_in[3];
  assign \dp/cache_in_mem_int[2]  = dcache_data_in[2];
  assign \dp/cache_in_mem_int[1]  = dcache_data_in[1];
  assign \dp/cache_in_mem_int[0]  = dcache_data_in[0];
  assign dcache_address[31] = \dp/mul_feedback_exe_mem_int[31] ;
  assign dcache_address[30] = \dp/mul_feedback_exe_mem_int[30] ;
  assign dcache_address[29] = \dp/mul_feedback_exe_mem_int[29] ;
  assign dcache_address[28] = \dp/mul_feedback_exe_mem_int[28] ;
  assign dcache_address[27] = \dp/mul_feedback_exe_mem_int[27] ;
  assign dcache_address[26] = \dp/mul_feedback_exe_mem_int[26] ;
  assign dcache_address[25] = \dp/mul_feedback_exe_mem_int[25] ;
  assign dcache_address[24] = \dp/mul_feedback_exe_mem_int[24] ;
  assign dcache_address[23] = \dp/mul_feedback_exe_mem_int[23] ;
  assign dcache_address[22] = \dp/mul_feedback_exe_mem_int[22] ;
  assign dcache_address[21] = \dp/mul_feedback_exe_mem_int[21] ;
  assign dcache_address[20] = \dp/mul_feedback_exe_mem_int[20] ;
  assign dcache_address[19] = \dp/mul_feedback_exe_mem_int[19] ;
  assign dcache_address[18] = \dp/mul_feedback_exe_mem_int[18] ;
  assign dcache_address[17] = \dp/mul_feedback_exe_mem_int[17] ;
  assign dcache_address[16] = \dp/mul_feedback_exe_mem_int[16] ;
  assign dcache_address[15] = \dp/mul_feedback_exe_mem_int[15] ;
  assign dcache_address[14] = \dp/mul_feedback_exe_mem_int[14] ;
  assign dcache_address[13] = \dp/mul_feedback_exe_mem_int[13] ;
  assign dcache_address[12] = \dp/mul_feedback_exe_mem_int[12] ;
  assign dcache_address[11] = \dp/mul_feedback_exe_mem_int[11] ;
  assign dcache_address[10] = \dp/mul_feedback_exe_mem_int[10] ;
  assign dcache_address[9] = \dp/mul_feedback_exe_mem_int[9] ;
  assign dcache_address[8] = \dp/mul_feedback_exe_mem_int[8] ;
  assign dcache_address[7] = \dp/mul_feedback_exe_mem_int[7] ;
  assign dcache_address[6] = \dp/mul_feedback_exe_mem_int[6] ;
  assign dcache_address[5] = \dp/mul_feedback_exe_mem_int[5] ;
  assign dcache_address[4] = \dp/mul_feedback_exe_mem_int[4] ;
  assign dcache_address[3] = \dp/mul_feedback_exe_mem_int[3] ;
  assign dcache_address[2] = \dp/mul_feedback_exe_mem_int[2] ;
  assign dcache_address[1] = \dp/mul_feedback_exe_mem_int[1] ;
  assign dcache_address[0] = \dp/mul_feedback_exe_mem_int[0] ;
  assign \dp/ifs/pc_btb[29]  = btb_cache_data_out_read[29];
  assign \dp/ifs/pc_btb[28]  = btb_cache_data_out_read[28];
  assign \dp/ifs/pc_btb[27]  = btb_cache_data_out_read[27];
  assign \dp/ifs/pc_btb[26]  = btb_cache_data_out_read[26];
  assign \dp/ifs/pc_btb[25]  = btb_cache_data_out_read[25];
  assign \dp/ifs/pc_btb[24]  = btb_cache_data_out_read[24];
  assign \dp/ifs/pc_btb[23]  = btb_cache_data_out_read[23];
  assign \dp/ifs/pc_btb[22]  = btb_cache_data_out_read[22];
  assign \dp/ifs/pc_btb[21]  = btb_cache_data_out_read[21];
  assign \dp/ifs/pc_btb[20]  = btb_cache_data_out_read[20];
  assign \dp/ifs/pc_btb[19]  = btb_cache_data_out_read[19];
  assign \dp/ifs/pc_btb[18]  = btb_cache_data_out_read[18];
  assign \dp/ifs/pc_btb[17]  = btb_cache_data_out_read[17];
  assign \dp/ifs/pc_btb[16]  = btb_cache_data_out_read[16];
  assign \dp/ifs/pc_btb[15]  = btb_cache_data_out_read[15];
  assign \dp/ifs/pc_btb[14]  = btb_cache_data_out_read[14];
  assign \dp/ifs/pc_btb[13]  = btb_cache_data_out_read[13];
  assign \dp/ifs/pc_btb[12]  = btb_cache_data_out_read[12];
  assign \dp/ifs/pc_btb[11]  = btb_cache_data_out_read[11];
  assign \dp/ifs/pc_btb[10]  = btb_cache_data_out_read[10];
  assign \dp/ifs/pc_btb[9]  = btb_cache_data_out_read[9];
  assign \dp/ifs/pc_btb[8]  = btb_cache_data_out_read[8];
  assign \dp/ifs/pc_btb[7]  = btb_cache_data_out_read[7];
  assign \dp/ifs/pc_btb[6]  = btb_cache_data_out_read[6];
  assign \dp/ifs/pc_btb[5]  = btb_cache_data_out_read[5];
  assign \dp/ifs/pc_btb[4]  = btb_cache_data_out_read[4];
  assign \dp/ifs/pc_btb[3]  = btb_cache_data_out_read[3];
  assign \dp/ifs/pc_btb[2]  = btb_cache_data_out_read[2];
  assign \dp/ifs/pc_btb[1]  = btb_cache_data_out_read[1];
  assign \dp/ifs/pc_btb[0]  = btb_cache_data_out_read[0];

  rf_N32 \dp/ids/reg_file  ( .clk(clk), .rst(rst_mem_wb_regs), .rp1_addr(rs_id), .rp2_addr(rt_id), .wp_addr({rd[4], n7535, rd[2:0]}), .wp_en(wp_en), .wp(
        wp_data), .rp1({\dp/ids/rp1[31] , \dp/ids/rp1[30] , \dp/ids/rp1[29] , 
        \dp/ids/rp1[28] , \dp/ids/rp1[27] , \dp/ids/rp1[26] , \dp/ids/rp1[25] , 
        \dp/ids/rp1[24] , \dp/ids/rp1[23] , \dp/ids/rp1[22] , \dp/ids/rp1[21] , 
        \dp/ids/rp1[20] , \dp/ids/rp1[19] , \dp/ids/rp1[18] , \dp/ids/rp1[17] , 
        \dp/ids/rp1[16] , \dp/ids/rp1[15] , \dp/ids/rp1[14] , \dp/ids/rp1[13] , 
        \dp/ids/rp1[12] , \dp/ids/rp1[11] , \dp/ids/rp1[10] , \dp/ids/rp1[9] , 
        \dp/ids/rp1[8] , \dp/ids/rp1[7] , \dp/ids/rp1[6] , \dp/ids/rp1[5] , 
        \dp/ids/rp1[4] , \dp/ids/rp1[3] , \dp/ids/rp1[2] , \dp/ids/rp1[1] , 
        \dp/ids/rp1[0] }), .rp2({\dp/ids/rp2[31] , \dp/ids/rp2[30] , 
        \dp/ids/rp2[29] , \dp/ids/rp2[28] , \dp/ids/rp2[27] , \dp/ids/rp2[26] , 
        \dp/ids/rp2[25] , \dp/ids/rp2[24] , \dp/ids/rp2[23] , \dp/ids/rp2[22] , 
        \dp/ids/rp2[21] , \dp/ids/rp2[20] , \dp/ids/rp2[19] , \dp/ids/rp2[18] , 
        \dp/ids/rp2[17] , \dp/ids/rp2[16] , \dp/ids/rp2[15] , \dp/ids/rp2[14] , 
        \dp/ids/rp2[13] , \dp/ids/rp2[12] , \dp/ids/rp2[11] , \dp/ids/rp2[10] , 
        \dp/ids/rp2[9] , \dp/ids/rp2[8] , \dp/ids/rp2[7] , \dp/ids/rp2[6] , 
        \dp/ids/rp2[5] , \dp/ids/rp2[4] , \dp/ids/rp2[3] , \dp/ids/rp2[2] , 
        \dp/ids/rp2[1] , \dp/ids/rp2[0] }), .rp1_out_sel(rp1_out_sel_id), 
        .rp2_out_sel(rp2_out_sel_id), .hilo_wr_en(hilo_wr_en), .lo_in({
        \dp/alu_out_low_mem_wb_int[31] , \dp/alu_out_low_mem_wb_int[30] , 
        \dp/alu_out_low_mem_wb_int[29] , \dp/alu_out_low_mem_wb_int[28] , 
        \dp/alu_out_low_mem_wb_int[27] , \dp/alu_out_low_mem_wb_int[26] , 
        \dp/alu_out_low_mem_wb_int[25] , \dp/alu_out_low_mem_wb_int[24] , 
        \dp/alu_out_low_mem_wb_int[23] , \dp/alu_out_low_mem_wb_int[22] , 
        \dp/alu_out_low_mem_wb_int[21] , \dp/alu_out_low_mem_wb_int[20] , 
        \dp/alu_out_low_mem_wb_int[19] , \dp/alu_out_low_mem_wb_int[18] , 
        \dp/alu_out_low_mem_wb_int[17] , \dp/alu_out_low_mem_wb_int[16] , 
        \dp/alu_out_low_mem_wb_int[15] , \dp/alu_out_low_mem_wb_int[14] , 
        \dp/alu_out_low_mem_wb_int[13] , \dp/alu_out_low_mem_wb_int[12] , 
        \dp/alu_out_low_mem_wb_int[11] , \dp/alu_out_low_mem_wb_int[10] , 
        \dp/alu_out_low_mem_wb_int[9] , \dp/alu_out_low_mem_wb_int[8] , 
        \dp/alu_out_low_mem_wb_int[7] , \dp/alu_out_low_mem_wb_int[6] , 
        \dp/alu_out_low_mem_wb_int[5] , \dp/alu_out_low_mem_wb_int[4] , 
        \dp/alu_out_low_mem_wb_int[3] , \dp/alu_out_low_mem_wb_int[2] , 
        \dp/alu_out_low_mem_wb_int[1] , \dp/alu_out_low_mem_wb_int[0] }), 
        .hi_in(wp_alu_data_high) );
  shifter_t2 \dp/exs/alu_unit/shifter  ( .data_in({\dp/exs/a_shift_int[31] , 
        \dp/exs/a_shift_int[30] , \dp/exs/a_shift_int[29] , 
        \dp/exs/a_shift_int[28] , \dp/exs/a_shift_int[27] , 
        \dp/exs/a_shift_int[26] , \dp/exs/a_shift_int[25] , 
        \dp/exs/a_shift_int[24] , \dp/exs/a_shift_int[23] , 
        \dp/exs/a_shift_int[22] , \dp/exs/a_shift_int[21] , 
        \dp/exs/a_shift_int[20] , \dp/exs/a_shift_int[19] , 
        \dp/exs/a_shift_int[18] , \dp/exs/a_shift_int[17] , 
        \dp/exs/a_shift_int[16] , \dp/exs/a_shift_int[15] , 
        \dp/exs/a_shift_int[14] , \dp/exs/a_shift_int[13] , 
        \dp/exs/a_shift_int[12] , \dp/exs/a_shift_int[11] , 
        \dp/exs/a_shift_int[10] , \dp/exs/a_shift_int[9] , 
        \dp/exs/a_shift_int[8] , \dp/exs/a_shift_int[7] , 
        \dp/exs/a_shift_int[6] , \dp/exs/a_shift_int[5] , 
        \dp/exs/a_shift_int[4] , \dp/exs/a_shift_int[3] , 
        \dp/exs/a_shift_int[2] , \dp/exs/a_shift_int[1] , 
        \dp/exs/a_shift_int[0] }), .shift({n110, n103, n99, n95, n92}), 
        .shift_type({1'b0, shift_type_exe[2:0]}), .data_out({
        \dp/exs/alu_unit/shifter_out[31] , \dp/exs/alu_unit/shifter_out[30] , 
        \dp/exs/alu_unit/shifter_out[29] , \dp/exs/alu_unit/shifter_out[28] , 
        \dp/exs/alu_unit/shifter_out[27] , \dp/exs/alu_unit/shifter_out[26] , 
        \dp/exs/alu_unit/shifter_out[25] , \dp/exs/alu_unit/shifter_out[24] , 
        \dp/exs/alu_unit/shifter_out[23] , \dp/exs/alu_unit/shifter_out[22] , 
        \dp/exs/alu_unit/shifter_out[21] , \dp/exs/alu_unit/shifter_out[20] , 
        \dp/exs/alu_unit/shifter_out[19] , \dp/exs/alu_unit/shifter_out[18] , 
        \dp/exs/alu_unit/shifter_out[17] , \dp/exs/alu_unit/shifter_out[16] , 
        \dp/exs/alu_unit/shifter_out[15] , \dp/exs/alu_unit/shifter_out[14] , 
        \dp/exs/alu_unit/shifter_out[13] , \dp/exs/alu_unit/shifter_out[12] , 
        \dp/exs/alu_unit/shifter_out[11] , \dp/exs/alu_unit/shifter_out[10] , 
        \dp/exs/alu_unit/shifter_out[9] , \dp/exs/alu_unit/shifter_out[8] , 
        \dp/exs/alu_unit/shifter_out[7] , \dp/exs/alu_unit/shifter_out[6] , 
        \dp/exs/alu_unit/shifter_out[5] , \dp/exs/alu_unit/shifter_out[4] , 
        \dp/exs/alu_unit/shifter_out[3] , \dp/exs/alu_unit/shifter_out[2] , 
        \dp/exs/alu_unit/shifter_out[1] , \dp/exs/alu_unit/shifter_out[0] })
         );
  a_generator \dp/exs/alu_unit/mult/a_gen  ( .a_in({1'b0, 1'b0, 
        \dp/a_mult_id_exe_int[61] , \dp/a_mult_id_exe_int[60] , 
        \dp/a_mult_id_exe_int[59] , \dp/a_mult_id_exe_int[58] , 
        \dp/a_mult_id_exe_int[57] , \dp/a_mult_id_exe_int[56] , 
        \dp/a_mult_id_exe_int[55] , \dp/a_mult_id_exe_int[54] , 
        \dp/a_mult_id_exe_int[53] , \dp/a_mult_id_exe_int[52] , 
        \dp/a_mult_id_exe_int[51] , \dp/a_mult_id_exe_int[50] , 
        \dp/a_mult_id_exe_int[49] , \dp/a_mult_id_exe_int[48] , 
        \dp/a_mult_id_exe_int[47] , \dp/a_mult_id_exe_int[46] , 
        \dp/a_mult_id_exe_int[45] , \dp/a_mult_id_exe_int[44] , 
        \dp/a_mult_id_exe_int[43] , \dp/a_mult_id_exe_int[42] , 
        \dp/a_mult_id_exe_int[41] , \dp/a_mult_id_exe_int[40] , 
        \dp/a_mult_id_exe_int[39] , \dp/a_mult_id_exe_int[38] , 
        \dp/a_mult_id_exe_int[37] , \dp/a_mult_id_exe_int[36] , 
        \dp/a_mult_id_exe_int[35] , \dp/a_mult_id_exe_int[34] , 
        \dp/a_mult_id_exe_int[33] , \dp/a_mult_id_exe_int[32] , 
        \dp/a_mult_id_exe_int[31] , \dp/a_mult_id_exe_int[30] , 
        \dp/a_mult_id_exe_int[29] , \dp/a_mult_id_exe_int[28] , 
        \dp/a_mult_id_exe_int[27] , \dp/a_mult_id_exe_int[26] , 
        \dp/a_mult_id_exe_int[25] , \dp/a_mult_id_exe_int[24] , 
        \dp/a_mult_id_exe_int[23] , \dp/a_mult_id_exe_int[22] , 
        \dp/a_mult_id_exe_int[21] , \dp/a_mult_id_exe_int[20] , 
        \dp/a_mult_id_exe_int[19] , \dp/a_mult_id_exe_int[18] , 
        \dp/a_mult_id_exe_int[17] , \dp/a_mult_id_exe_int[16] , 
        \dp/a_mult_id_exe_int[15] , \dp/a_mult_id_exe_int[14] , 
        \dp/a_mult_id_exe_int[13] , \dp/a_mult_id_exe_int[12] , 
        \dp/a_mult_id_exe_int[11] , \dp/a_mult_id_exe_int[10] , 
        \dp/a_mult_id_exe_int[9] , \dp/a_mult_id_exe_int[8] , 
        \dp/a_mult_id_exe_int[7] , \dp/a_mult_id_exe_int[6] , 
        \dp/a_mult_id_exe_int[5] , \dp/a_mult_id_exe_int[4] , 
        \dp/a_mult_id_exe_int[3] , \dp/a_mult_id_exe_int[2] , 
        \dp/a_mult_id_exe_int[1] , \dp/a_mult_id_exe_int[0] }), .neg_a_in({
        1'b0, 1'b0, \dp/a_neg_mult_id_exe_int[61] , 
        \dp/a_neg_mult_id_exe_int[60] , \dp/a_neg_mult_id_exe_int[59] , 
        \dp/a_neg_mult_id_exe_int[58] , \dp/a_neg_mult_id_exe_int[57] , 
        \dp/a_neg_mult_id_exe_int[56] , \dp/a_neg_mult_id_exe_int[55] , 
        \dp/a_neg_mult_id_exe_int[54] , \dp/a_neg_mult_id_exe_int[53] , 
        \dp/a_neg_mult_id_exe_int[52] , \dp/a_neg_mult_id_exe_int[51] , 
        \dp/a_neg_mult_id_exe_int[50] , \dp/a_neg_mult_id_exe_int[49] , 
        \dp/a_neg_mult_id_exe_int[48] , \dp/a_neg_mult_id_exe_int[47] , 
        \dp/a_neg_mult_id_exe_int[46] , \dp/a_neg_mult_id_exe_int[45] , 
        \dp/a_neg_mult_id_exe_int[44] , \dp/a_neg_mult_id_exe_int[43] , 
        \dp/a_neg_mult_id_exe_int[42] , \dp/a_neg_mult_id_exe_int[41] , 
        \dp/a_neg_mult_id_exe_int[40] , \dp/a_neg_mult_id_exe_int[39] , 
        \dp/a_neg_mult_id_exe_int[38] , \dp/a_neg_mult_id_exe_int[37] , 
        \dp/a_neg_mult_id_exe_int[36] , \dp/a_neg_mult_id_exe_int[35] , 
        \dp/a_neg_mult_id_exe_int[34] , \dp/a_neg_mult_id_exe_int[33] , 
        \dp/a_neg_mult_id_exe_int[32] , \dp/a_neg_mult_id_exe_int[31] , 
        \dp/a_neg_mult_id_exe_int[30] , \dp/a_neg_mult_id_exe_int[29] , 
        \dp/a_neg_mult_id_exe_int[28] , \dp/a_neg_mult_id_exe_int[27] , 
        \dp/a_neg_mult_id_exe_int[26] , \dp/a_neg_mult_id_exe_int[25] , 
        \dp/a_neg_mult_id_exe_int[24] , \dp/a_neg_mult_id_exe_int[23] , 
        \dp/a_neg_mult_id_exe_int[22] , \dp/a_neg_mult_id_exe_int[21] , 
        \dp/a_neg_mult_id_exe_int[20] , \dp/a_neg_mult_id_exe_int[19] , 
        \dp/a_neg_mult_id_exe_int[18] , \dp/a_neg_mult_id_exe_int[17] , 
        \dp/a_neg_mult_id_exe_int[16] , \dp/a_neg_mult_id_exe_int[15] , 
        \dp/a_neg_mult_id_exe_int[14] , \dp/a_neg_mult_id_exe_int[13] , 
        \dp/a_neg_mult_id_exe_int[12] , \dp/a_neg_mult_id_exe_int[11] , 
        \dp/a_neg_mult_id_exe_int[10] , \dp/a_neg_mult_id_exe_int[9] , 
        \dp/a_neg_mult_id_exe_int[8] , \dp/a_neg_mult_id_exe_int[7] , 
        \dp/a_neg_mult_id_exe_int[6] , \dp/a_neg_mult_id_exe_int[5] , 
        \dp/a_neg_mult_id_exe_int[4] , \dp/a_neg_mult_id_exe_int[3] , 
        \dp/a_neg_mult_id_exe_int[2] , \dp/a_neg_mult_id_exe_int[1] , 
        \dp/a_neg_mult_id_exe_int[0] }), .sel({it_exe[3:1], n5159}), .a({
        \dp/exs/alu_unit/mult/a_shiftn[63] , 
        \dp/exs/alu_unit/mult/a_shiftn[62] , 
        \dp/exs/alu_unit/mult/a_shiftn[61] , 
        \dp/exs/alu_unit/mult/a_shiftn[60] , 
        \dp/exs/alu_unit/mult/a_shiftn[59] , 
        \dp/exs/alu_unit/mult/a_shiftn[58] , 
        \dp/exs/alu_unit/mult/a_shiftn[57] , 
        \dp/exs/alu_unit/mult/a_shiftn[56] , 
        \dp/exs/alu_unit/mult/a_shiftn[55] , 
        \dp/exs/alu_unit/mult/a_shiftn[54] , 
        \dp/exs/alu_unit/mult/a_shiftn[53] , 
        \dp/exs/alu_unit/mult/a_shiftn[52] , 
        \dp/exs/alu_unit/mult/a_shiftn[51] , 
        \dp/exs/alu_unit/mult/a_shiftn[50] , 
        \dp/exs/alu_unit/mult/a_shiftn[49] , 
        \dp/exs/alu_unit/mult/a_shiftn[48] , 
        \dp/exs/alu_unit/mult/a_shiftn[47] , 
        \dp/exs/alu_unit/mult/a_shiftn[46] , 
        \dp/exs/alu_unit/mult/a_shiftn[45] , 
        \dp/exs/alu_unit/mult/a_shiftn[44] , 
        \dp/exs/alu_unit/mult/a_shiftn[43] , 
        \dp/exs/alu_unit/mult/a_shiftn[42] , 
        \dp/exs/alu_unit/mult/a_shiftn[41] , 
        \dp/exs/alu_unit/mult/a_shiftn[40] , 
        \dp/exs/alu_unit/mult/a_shiftn[39] , 
        \dp/exs/alu_unit/mult/a_shiftn[38] , 
        \dp/exs/alu_unit/mult/a_shiftn[37] , 
        \dp/exs/alu_unit/mult/a_shiftn[36] , 
        \dp/exs/alu_unit/mult/a_shiftn[35] , 
        \dp/exs/alu_unit/mult/a_shiftn[34] , 
        \dp/exs/alu_unit/mult/a_shiftn[33] , 
        \dp/exs/alu_unit/mult/a_shiftn[32] , 
        \dp/exs/alu_unit/mult/a_shiftn[31] , 
        \dp/exs/alu_unit/mult/a_shiftn[30] , 
        \dp/exs/alu_unit/mult/a_shiftn[29] , 
        \dp/exs/alu_unit/mult/a_shiftn[28] , 
        \dp/exs/alu_unit/mult/a_shiftn[27] , 
        \dp/exs/alu_unit/mult/a_shiftn[26] , 
        \dp/exs/alu_unit/mult/a_shiftn[25] , 
        \dp/exs/alu_unit/mult/a_shiftn[24] , 
        \dp/exs/alu_unit/mult/a_shiftn[23] , 
        \dp/exs/alu_unit/mult/a_shiftn[22] , 
        \dp/exs/alu_unit/mult/a_shiftn[21] , 
        \dp/exs/alu_unit/mult/a_shiftn[20] , 
        \dp/exs/alu_unit/mult/a_shiftn[19] , 
        \dp/exs/alu_unit/mult/a_shiftn[18] , 
        \dp/exs/alu_unit/mult/a_shiftn[17] , 
        \dp/exs/alu_unit/mult/a_shiftn[16] , 
        \dp/exs/alu_unit/mult/a_shiftn[15] , 
        \dp/exs/alu_unit/mult/a_shiftn[14] , 
        \dp/exs/alu_unit/mult/a_shiftn[13] , 
        \dp/exs/alu_unit/mult/a_shiftn[12] , SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        \dp/exs/alu_unit/mult/a_shiftn[2] , SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10}), .neg_a({
        \dp/exs/alu_unit/mult/neg_a_shiftn[63] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[62] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[61] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[60] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[59] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[58] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[57] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[56] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[55] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[54] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[53] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[52] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[51] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[50] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[49] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[48] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[47] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[46] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[45] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[44] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[43] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[42] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[41] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[40] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[39] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[38] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[37] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[36] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[35] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[34] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[33] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[32] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[31] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[30] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[29] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[28] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[27] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[26] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[25] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[24] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[23] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[22] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[21] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[20] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[19] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[18] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[17] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[16] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[15] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[14] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[13] , 
        \dp/exs/alu_unit/mult/neg_a_shiftn[12] , SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        \dp/exs/alu_unit/mult/neg_a_shiftn[2] , SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21}), .ax2({SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, SYNOPSYS_UNCONNECTED__32, 
        SYNOPSYS_UNCONNECTED__33, SYNOPSYS_UNCONNECTED__34, 
        SYNOPSYS_UNCONNECTED__35, SYNOPSYS_UNCONNECTED__36, 
        SYNOPSYS_UNCONNECTED__37, SYNOPSYS_UNCONNECTED__38, 
        SYNOPSYS_UNCONNECTED__39, SYNOPSYS_UNCONNECTED__40, 
        SYNOPSYS_UNCONNECTED__41, SYNOPSYS_UNCONNECTED__42, 
        SYNOPSYS_UNCONNECTED__43, SYNOPSYS_UNCONNECTED__44, 
        SYNOPSYS_UNCONNECTED__45, SYNOPSYS_UNCONNECTED__46, 
        SYNOPSYS_UNCONNECTED__47, SYNOPSYS_UNCONNECTED__48, 
        SYNOPSYS_UNCONNECTED__49, SYNOPSYS_UNCONNECTED__50, 
        SYNOPSYS_UNCONNECTED__51, SYNOPSYS_UNCONNECTED__52, 
        SYNOPSYS_UNCONNECTED__53, SYNOPSYS_UNCONNECTED__54, 
        SYNOPSYS_UNCONNECTED__55, SYNOPSYS_UNCONNECTED__56, 
        SYNOPSYS_UNCONNECTED__57, SYNOPSYS_UNCONNECTED__58, 
        SYNOPSYS_UNCONNECTED__59, SYNOPSYS_UNCONNECTED__60, 
        SYNOPSYS_UNCONNECTED__61, SYNOPSYS_UNCONNECTED__62, 
        SYNOPSYS_UNCONNECTED__63, SYNOPSYS_UNCONNECTED__64, 
        SYNOPSYS_UNCONNECTED__65, SYNOPSYS_UNCONNECTED__66, 
        SYNOPSYS_UNCONNECTED__67, SYNOPSYS_UNCONNECTED__68, 
        SYNOPSYS_UNCONNECTED__69, SYNOPSYS_UNCONNECTED__70, 
        SYNOPSYS_UNCONNECTED__71, SYNOPSYS_UNCONNECTED__72, 
        \dp/exs/alu_unit/mult/ax2_shiftn[12] , 
        \dp/exs/alu_unit/mult/ax2_shiftn[11] , 
        \dp/exs/alu_unit/mult/ax2_shiftn[10] , 
        \dp/exs/alu_unit/mult/ax2_shiftn[9] , 
        \dp/exs/alu_unit/mult/ax2_shiftn[8] , 
        \dp/exs/alu_unit/mult/ax2_shiftn[7] , 
        \dp/exs/alu_unit/mult/ax2_shiftn[6] , 
        \dp/exs/alu_unit/mult/ax2_shiftn[5] , 
        \dp/exs/alu_unit/mult/ax2_shiftn[4] , SYNOPSYS_UNCONNECTED__73, 
        SYNOPSYS_UNCONNECTED__74, SYNOPSYS_UNCONNECTED__75, 
        SYNOPSYS_UNCONNECTED__76}), .neg_ax2({SYNOPSYS_UNCONNECTED__77, 
        SYNOPSYS_UNCONNECTED__78, SYNOPSYS_UNCONNECTED__79, 
        SYNOPSYS_UNCONNECTED__80, SYNOPSYS_UNCONNECTED__81, 
        SYNOPSYS_UNCONNECTED__82, SYNOPSYS_UNCONNECTED__83, 
        SYNOPSYS_UNCONNECTED__84, SYNOPSYS_UNCONNECTED__85, 
        SYNOPSYS_UNCONNECTED__86, SYNOPSYS_UNCONNECTED__87, 
        SYNOPSYS_UNCONNECTED__88, SYNOPSYS_UNCONNECTED__89, 
        SYNOPSYS_UNCONNECTED__90, SYNOPSYS_UNCONNECTED__91, 
        SYNOPSYS_UNCONNECTED__92, SYNOPSYS_UNCONNECTED__93, 
        SYNOPSYS_UNCONNECTED__94, SYNOPSYS_UNCONNECTED__95, 
        SYNOPSYS_UNCONNECTED__96, SYNOPSYS_UNCONNECTED__97, 
        SYNOPSYS_UNCONNECTED__98, SYNOPSYS_UNCONNECTED__99, 
        SYNOPSYS_UNCONNECTED__100, SYNOPSYS_UNCONNECTED__101, 
        SYNOPSYS_UNCONNECTED__102, SYNOPSYS_UNCONNECTED__103, 
        SYNOPSYS_UNCONNECTED__104, SYNOPSYS_UNCONNECTED__105, 
        SYNOPSYS_UNCONNECTED__106, SYNOPSYS_UNCONNECTED__107, 
        SYNOPSYS_UNCONNECTED__108, SYNOPSYS_UNCONNECTED__109, 
        SYNOPSYS_UNCONNECTED__110, SYNOPSYS_UNCONNECTED__111, 
        SYNOPSYS_UNCONNECTED__112, SYNOPSYS_UNCONNECTED__113, 
        SYNOPSYS_UNCONNECTED__114, SYNOPSYS_UNCONNECTED__115, 
        SYNOPSYS_UNCONNECTED__116, SYNOPSYS_UNCONNECTED__117, 
        SYNOPSYS_UNCONNECTED__118, SYNOPSYS_UNCONNECTED__119, 
        SYNOPSYS_UNCONNECTED__120, SYNOPSYS_UNCONNECTED__121, 
        SYNOPSYS_UNCONNECTED__122, SYNOPSYS_UNCONNECTED__123, 
        SYNOPSYS_UNCONNECTED__124, SYNOPSYS_UNCONNECTED__125, 
        SYNOPSYS_UNCONNECTED__126, SYNOPSYS_UNCONNECTED__127, 
        \dp/exs/alu_unit/mult/neg_ax2_shiftn[12] , 
        \dp/exs/alu_unit/mult/neg_ax2_shiftn[11] , 
        \dp/exs/alu_unit/mult/neg_ax2_shiftn[10] , 
        \dp/exs/alu_unit/mult/neg_ax2_shiftn[9] , 
        \dp/exs/alu_unit/mult/neg_ax2_shiftn[8] , 
        \dp/exs/alu_unit/mult/neg_ax2_shiftn[7] , 
        \dp/exs/alu_unit/mult/neg_ax2_shiftn[6] , 
        \dp/exs/alu_unit/mult/neg_ax2_shiftn[5] , 
        \dp/exs/alu_unit/mult/neg_ax2_shiftn[4] , SYNOPSYS_UNCONNECTED__128, 
        SYNOPSYS_UNCONNECTED__129, SYNOPSYS_UNCONNECTED__130, 
        SYNOPSYS_UNCONNECTED__131}) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[15]  ( .D(n3131), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[15] ), .QN(n4538) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[14]  ( .D(n3132), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[14] ), .QN(n4529) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[13]  ( .D(n3133), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[13] ), .QN(n4528) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[12]  ( .D(n3134), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[12] ), .QN(n4527) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[11]  ( .D(n3135), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[11] ), .QN(n4526) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[10]  ( .D(n3136), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[10] ), .QN(n4525) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[9]  ( .D(n3137), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[9] ), .QN(n4524) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[8]  ( .D(n3138), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[8] ), .QN(n4523) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[31]  ( .D(n3115), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[31] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[30]  ( .D(n3116), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[30] ), .QN(n4277) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[29]  ( .D(n3117), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[29] ), .QN(n4278) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[28]  ( .D(n3118), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[28] ), .QN(n4279) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[27]  ( .D(n3119), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[27] ), .QN(n4280) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[26]  ( .D(n3120), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[26] ), .QN(n4281) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[25]  ( .D(n3121), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[25] ), .QN(n4282) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[24]  ( .D(n3122), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[24] ), .QN(n4283) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[23]  ( .D(n3123), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[23] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[22]  ( .D(n3124), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[22] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[21]  ( .D(n3125), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[21] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[20]  ( .D(n3126), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[20] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[19]  ( .D(n3127), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[19] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[18]  ( .D(n3128), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[18] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[17]  ( .D(n3129), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[17] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[16]  ( .D(n3130), .CK(clk), .Q(
        \dp/cache_data_mem_wb_int[16] ) );
  DFF_X1 \mc/currstate_reg[0]  ( .D(n3114), .CK(clk), .Q(\mc/currstate[0] ), 
        .QN(n4371) );
  DFF_X1 \mc/curr_cache_data_reg[31]  ( .D(n3073), .CK(clk), .Q(n4637), .QN(
        n330) );
  DFF_X1 \mc/curr_cache_data_reg[30]  ( .D(n3074), .CK(clk), .Q(n4636), .QN(
        n329) );
  DFF_X1 \mc/curr_cache_data_reg[29]  ( .D(n3075), .CK(clk), .Q(n4635), .QN(
        n328) );
  DFF_X1 \mc/curr_cache_data_reg[28]  ( .D(n3076), .CK(clk), .Q(n4634), .QN(
        n327) );
  DFF_X1 \mc/curr_cache_data_reg[27]  ( .D(n3077), .CK(clk), .Q(n4633), .QN(
        n326) );
  DFF_X1 \mc/curr_cache_data_reg[26]  ( .D(n3078), .CK(clk), .Q(n4632), .QN(
        n325) );
  DFF_X1 \mc/curr_cache_data_reg[25]  ( .D(n3079), .CK(clk), .Q(n4631), .QN(
        n324) );
  DFF_X1 \mc/curr_cache_data_reg[24]  ( .D(n3080), .CK(clk), .Q(n4630), .QN(
        n323) );
  DFF_X1 \mc/curr_cache_data_reg[23]  ( .D(n3081), .CK(clk), .Q(n4629), .QN(
        n322) );
  DFF_X1 \mc/curr_cache_data_reg[22]  ( .D(n3082), .CK(clk), .Q(n4628), .QN(
        n321) );
  DFF_X1 \mc/curr_cache_data_reg[21]  ( .D(n3083), .CK(clk), .Q(n4627), .QN(
        n320) );
  DFF_X1 \mc/curr_cache_data_reg[20]  ( .D(n3084), .CK(clk), .Q(n4626), .QN(
        n319) );
  DFF_X1 \mc/curr_cache_data_reg[19]  ( .D(n3085), .CK(clk), .Q(n4625), .QN(
        n318) );
  DFF_X1 \mc/curr_cache_data_reg[18]  ( .D(n3086), .CK(clk), .Q(n4624), .QN(
        n317) );
  DFF_X1 \mc/curr_cache_data_reg[17]  ( .D(n3087), .CK(clk), .Q(n4623), .QN(
        n316) );
  DFF_X1 \mc/curr_cache_data_reg[16]  ( .D(n3088), .CK(clk), .Q(n4622), .QN(
        n315) );
  DFF_X1 \mc/curr_cache_data_reg[15]  ( .D(n3089), .CK(clk), .Q(n4621), .QN(
        n314) );
  DFF_X1 \mc/curr_cache_data_reg[14]  ( .D(n3090), .CK(clk), .Q(n4620), .QN(
        n313) );
  DFF_X1 \mc/curr_cache_data_reg[13]  ( .D(n3091), .CK(clk), .Q(n4619), .QN(
        n312) );
  DFF_X1 \mc/curr_cache_data_reg[12]  ( .D(n3092), .CK(clk), .Q(n4618), .QN(
        n311) );
  DFF_X1 \mc/curr_cache_data_reg[11]  ( .D(n3093), .CK(clk), .Q(n4617), .QN(
        n310) );
  DFF_X1 \mc/curr_cache_data_reg[10]  ( .D(n3094), .CK(clk), .Q(n4616), .QN(
        n309) );
  DFF_X1 \mc/curr_cache_data_reg[9]  ( .D(n3095), .CK(clk), .Q(n4615), .QN(
        n308) );
  DFF_X1 \mc/curr_cache_data_reg[8]  ( .D(n3096), .CK(clk), .Q(n4614), .QN(
        n307) );
  DFF_X1 \mc/curr_cache_data_reg[7]  ( .D(n3097), .CK(clk), .Q(n4613), .QN(
        n306) );
  DFF_X1 \mc/curr_cache_data_reg[6]  ( .D(n3098), .CK(clk), .Q(n4612), .QN(
        n305) );
  DFF_X1 \mc/curr_cache_data_reg[5]  ( .D(n3099), .CK(clk), .Q(n4611), .QN(
        n304) );
  DFF_X1 \mc/curr_cache_data_reg[4]  ( .D(n3100), .CK(clk), .Q(n4610), .QN(
        n303) );
  DFF_X1 \mc/curr_cache_data_reg[3]  ( .D(n3101), .CK(clk), .Q(n4609), .QN(
        n302) );
  DFF_X1 \mc/curr_cache_data_reg[2]  ( .D(n3102), .CK(clk), .Q(n4608), .QN(
        n301) );
  DFF_X1 \mc/curr_cache_data_reg[1]  ( .D(n3103), .CK(clk), .Q(n4607), .QN(
        n300) );
  DFF_X1 \mc/curr_cache_data_reg[0]  ( .D(n3104), .CK(clk), .Q(n4606), .QN(
        n299) );
  DFF_X1 \mc/curr_evicted_address_reg[7]  ( .D(n3105), .CK(clk), .Q(n4645), 
        .QN(n295) );
  DFF_X1 \mc/curr_evicted_address_reg[6]  ( .D(n3106), .CK(clk), .Q(n4644), 
        .QN(n294) );
  DFF_X1 \mc/curr_evicted_address_reg[5]  ( .D(n3107), .CK(clk), .Q(n4643), 
        .QN(n293) );
  DFF_X1 \mc/curr_evicted_address_reg[4]  ( .D(n3108), .CK(clk), .Q(n4642), 
        .QN(n292) );
  DFF_X1 \mc/curr_evicted_address_reg[3]  ( .D(n3109), .CK(clk), .Q(n4641), 
        .QN(n291) );
  DFF_X1 \mc/curr_evicted_address_reg[2]  ( .D(n3110), .CK(clk), .Q(n4640), 
        .QN(n290) );
  DFF_X1 \mc/curr_evicted_address_reg[1]  ( .D(n3111), .CK(clk), .Q(n4639), 
        .QN(n289) );
  DFF_X1 \mc/curr_evicted_address_reg[0]  ( .D(n3112), .CK(clk), .Q(n4638), 
        .QN(n288) );
  DFF_X1 \mc/currstate_reg[1]  ( .D(n3113), .CK(clk), .Q(\mc/currstate[1] ), 
        .QN(n4266) );
  DFF_X1 \dp/id_exe_regs/rs_reg/q_reg[4]  ( .D(n3058), .CK(clk), .Q(rs_exe[4]), 
        .QN(n4500) );
  DFF_X1 \dp/id_exe_regs/rs_reg/q_reg[3]  ( .D(n3059), .CK(clk), .Q(rs_exe[3]), 
        .QN(n4490) );
  DFF_X1 \dp/id_exe_regs/rs_reg/q_reg[2]  ( .D(n3060), .CK(clk), .Q(rs_exe[2]), 
        .QN(n4499) );
  DFF_X1 \dp/id_exe_regs/rs_reg/q_reg[1]  ( .D(n3061), .CK(clk), .Q(rs_exe[1]), 
        .QN(n4489) );
  DFF_X1 \dp/id_exe_regs/rs_reg/q_reg[0]  ( .D(n3062), .CK(clk), .Q(rs_exe[0]), 
        .QN(n4498) );
  DFF_X1 \dp/id_exe_regs/rt_reg/q_reg[4]  ( .D(n3068), .CK(clk), .Q(rt_exe[4]), 
        .QN(n4497) );
  DFF_X1 \dp/id_exe_regs/rt_reg/q_reg[3]  ( .D(n3069), .CK(clk), .Q(rt_exe[3]), 
        .QN(n4496) );
  DFF_X1 \dp/id_exe_regs/rt_reg/q_reg[2]  ( .D(n3070), .CK(clk), .Q(rt_exe[2]), 
        .QN(n4495) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[17]  ( .D(n275), .CK(clk), .Q(rt_id[1]), 
        .QN(n4138) );
  DFF_X1 \dp/id_exe_regs/rt_reg/q_reg[1]  ( .D(n3071), .CK(clk), .Q(rt_exe[1]), 
        .QN(n4518) );
  DFF_X1 \dp/id_exe_regs/rt_reg/q_reg[0]  ( .D(n3072), .CK(clk), .Q(rt_exe[0]), 
        .QN(n4517) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[15]  ( .D(n1627), .CK(clk), .Q(n4368), 
        .QN(\dp/imm_id_int[15] ) );
  DFF_X1 \dp/id_exe_regs/rd_reg/q_reg[4]  ( .D(n3063), .CK(clk), .Q(
        rd_idexe[4]) );
  DFF_X1 \dp/ex_mem_regs/rd_reg/q_reg[4]  ( .D(n1600), .CK(clk), .Q(n4020), 
        .QN(rd_exemem[4]) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[15]  ( .D(n265), .CK(clk), .Q(
        \dp/imm_id_exe_int[15] ), .QN(n4070) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[23]  ( .D(n3050), .CK(clk), .Q(
        \dp/imm_id_exe_int[23] ), .QN(n3866) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[22]  ( .D(n3051), .CK(clk), .Q(
        \dp/imm_id_exe_int[22] ), .QN(n4220) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[21]  ( .D(n3052), .CK(clk), .Q(
        \dp/imm_id_exe_int[21] ), .QN(n4222) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[31]  ( .D(n3042), .CK(clk), .Q(
        \dp/imm_id_exe_int[31] ), .QN(n4503) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[30]  ( .D(n3043), .CK(clk), .Q(
        \dp/imm_id_exe_int[30] ), .QN(n4367) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[14]  ( .D(n1628), .CK(clk), .Q(n4364), 
        .QN(\dp/imm_id_int[14] ) );
  DFF_X1 \dp/id_exe_regs/rd_reg/q_reg[3]  ( .D(n3064), .CK(clk), .Q(
        rd_idexe[3]) );
  DFF_X1 \dp/ex_mem_regs/rd_reg/q_reg[3]  ( .D(n1603), .CK(clk), .Q(n4009), 
        .QN(rd_exemem[3]) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[14]  ( .D(n264), .CK(clk), .QN(n4118)
         );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[13]  ( .D(n1629), .CK(clk), .Q(n4363), 
        .QN(\dp/imm_id_int[13] ) );
  DFF_X1 \dp/id_exe_regs/rd_reg/q_reg[2]  ( .D(n3065), .CK(clk), .Q(
        rd_idexe[2]) );
  DFF_X1 \dp/ex_mem_regs/rd_reg/q_reg[2]  ( .D(n1604), .CK(clk), .Q(n4007), 
        .QN(rd_exemem[2]) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[13]  ( .D(n263), .CK(clk), .QN(n4119)
         );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[12]  ( .D(n1630), .CK(clk), .Q(n4362), 
        .QN(\dp/imm_id_int[12] ) );
  DFF_X1 \dp/id_exe_regs/rd_reg/q_reg[1]  ( .D(n3066), .CK(clk), .Q(
        rd_idexe[1]) );
  DFF_X1 \dp/ex_mem_regs/rd_reg/q_reg[1]  ( .D(n1605), .CK(clk), .QN(
        rd_exemem[1]) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[12]  ( .D(n262), .CK(clk), .QN(n4120)
         );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[11]  ( .D(n1631), .CK(clk), .Q(n4361), 
        .QN(\dp/imm_id_int[11] ) );
  DFF_X1 \dp/id_exe_regs/rd_reg/q_reg[0]  ( .D(n3067), .CK(clk), .Q(
        rd_idexe[0]), .QN(n4240) );
  DFF_X1 \dp/ex_mem_regs/rd_reg/q_reg[0]  ( .D(n1606), .CK(clk), .Q(n4018), 
        .QN(rd_exemem[0]) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[11]  ( .D(n261), .CK(clk), .QN(
        \intadd_2/A[8] ) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[10]  ( .D(n1632), .CK(clk), .Q(n4372), 
        .QN(\dp/imm_id_int[10] ) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[10]  ( .D(n260), .CK(clk), .QN(n4121)
         );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[9]  ( .D(n1633), .CK(clk), .Q(n4373), 
        .QN(\dp/imm_id_int[9] ) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[8]  ( .D(n1634), .CK(clk), .Q(n4374), 
        .QN(\dp/imm_id_int[8] ) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[8]  ( .D(n258), .CK(clk), .Q(
        \dp/imm_id_exe_int[8] ), .QN(n4098) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[7]  ( .D(n1635), .CK(clk), .Q(n4375), 
        .QN(\dp/imm_id_int[7] ) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[7]  ( .D(n257), .CK(clk), .Q(n4130), 
        .QN(\intadd_2/A[4] ) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[6]  ( .D(n1636), .CK(clk), .Q(n4376), 
        .QN(\dp/imm_id_int[6] ) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[6]  ( .D(n256), .CK(clk), .Q(
        \dp/imm_id_exe_int[6] ), .QN(n4099) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[5]  ( .D(n1637), .CK(clk), .Q(n4381), 
        .QN(\dp/imm_id_int[5] ) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[5]  ( .D(n255), .CK(clk), .Q(n4125), 
        .QN(\intadd_2/A[2] ) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[4]  ( .D(n1638), .CK(clk), .Q(n4447), 
        .QN(\dp/imm_id_int[4] ) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[4]  ( .D(n254), .CK(clk), .Q(
        \dp/imm_id_exe_int[4] ), .QN(n4100) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[3]  ( .D(n1639), .CK(clk), .Q(n4446), 
        .QN(\dp/imm_id_int[3] ) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[3]  ( .D(n253), .CK(clk), .QN(
        \intadd_2/A[0] ) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[2]  ( .D(n1640), .CK(clk), .Q(n4168), 
        .QN(\dp/imm_id_int[2] ) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[2]  ( .D(n252), .CK(clk), .Q(
        \dp/imm_id_exe_int[2] ), .QN(n4501) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[1]  ( .D(n1641), .CK(clk), .Q(n4476), 
        .QN(\dp/imm_id_int[1] ) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[0]  ( .D(n1642), .CK(clk), .Q(n4477), 
        .QN(\dp/imm_id_int[0] ) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[29]  ( .D(n3011), .CK(clk), .Q(n4384), 
        .QN(n389) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[31]  ( .D(n2979), .CK(clk), .Q(
        \dp/npc_id_exe_int[31] ), .QN(n4483) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[28]  ( .D(n3012), .CK(clk), .Q(n4408), 
        .QN(n388) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[30]  ( .D(n2980), .CK(clk), .Q(n4140), 
        .QN(n4519) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[27]  ( .D(n3013), .CK(clk), .Q(n4415), 
        .QN(n387) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[29]  ( .D(n2981), .CK(clk), .QN(n4536)
         );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[26]  ( .D(n3014), .CK(clk), .Q(n4416), 
        .QN(n386) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[28]  ( .D(n2982), .CK(clk), .Q(
        \dp/npc_id_exe_int[28] ), .QN(n4148) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[25]  ( .D(n3015), .CK(clk), .Q(n4417), 
        .QN(n385) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[27]  ( .D(n2983), .CK(clk), .QN(n4520)
         );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[24]  ( .D(n3016), .CK(clk), .Q(n4418), 
        .QN(n384) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[26]  ( .D(n2984), .CK(clk), .Q(
        \dp/npc_id_exe_int[26] ), .QN(n4147) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[23]  ( .D(n3017), .CK(clk), .Q(n4409), 
        .QN(n383) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[25]  ( .D(n2985), .CK(clk), .Q(
        \dp/npc_id_exe_int[25] ), .QN(n4137) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[22]  ( .D(n3018), .CK(clk), .Q(n4419), 
        .QN(n382) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[24]  ( .D(n2986), .CK(clk), .Q(
        \dp/npc_id_exe_int[24] ), .QN(n4356) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[21]  ( .D(n3019), .CK(clk), .Q(n4420), 
        .QN(n381) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[23]  ( .D(n2987), .CK(clk), .Q(
        \dp/npc_id_exe_int[23] ), .QN(\intadd_2/B[20] ) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[20]  ( .D(n3020), .CK(clk), .Q(n4443), 
        .QN(n380) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[22]  ( .D(n2988), .CK(clk), .Q(
        \dp/npc_id_exe_int[22] ), .QN(n4103) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[19]  ( .D(n3021), .CK(clk), .Q(n4421), 
        .QN(n379) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[21]  ( .D(n2989), .CK(clk), .Q(
        \dp/npc_id_exe_int[21] ), .QN(n4101) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[18]  ( .D(n3022), .CK(clk), .Q(n4422), 
        .QN(n378) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[20]  ( .D(n2990), .CK(clk), .Q(
        \dp/npc_id_exe_int[20] ), .QN(n4114) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[17]  ( .D(n3023), .CK(clk), .Q(n4423), 
        .QN(n377) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[19]  ( .D(n2991), .CK(clk), .QN(n4110)
         );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[16]  ( .D(n3024), .CK(clk), .Q(n4424), 
        .QN(n376) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[18]  ( .D(n2992), .CK(clk), .Q(
        \dp/npc_id_exe_int[18] ), .QN(n4113) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[15]  ( .D(n3025), .CK(clk), .Q(n4410), 
        .QN(n375) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[17]  ( .D(n2993), .CK(clk), .Q(
        \dp/npc_id_exe_int[17] ), .QN(\intadd_2/B[14] ) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[14]  ( .D(n3026), .CK(clk), .Q(n4411), 
        .QN(n374) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[16]  ( .D(n2994), .CK(clk), .Q(
        \dp/npc_id_exe_int[16] ), .QN(n4102) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[13]  ( .D(n3027), .CK(clk), .Q(n4425), 
        .QN(n373) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[15]  ( .D(n2995), .CK(clk), .Q(n4116), 
        .QN(n4207) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[12]  ( .D(n3028), .CK(clk), .Q(n4426), 
        .QN(n372) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[14]  ( .D(n2996), .CK(clk), .Q(
        \dp/npc_id_exe_int[14] ), .QN(n4235) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[11]  ( .D(n3029), .CK(clk), .Q(n4427), 
        .QN(n371) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[13]  ( .D(n2997), .CK(clk), .QN(n4226)
         );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[10]  ( .D(n3030), .CK(clk), .Q(n4428), 
        .QN(n370) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[12]  ( .D(n2998), .CK(clk), .Q(
        \dp/npc_id_exe_int[12] ), .QN(n4234) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[9]  ( .D(n3031), .CK(clk), .Q(n4429), 
        .QN(n369) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[11]  ( .D(n2999), .CK(clk), .QN(n4218)
         );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[8]  ( .D(n3032), .CK(clk), .Q(n4430), 
        .QN(n368) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[10]  ( .D(n3000), .CK(clk), .Q(
        \dp/npc_id_exe_int[10] ), .QN(n4233) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[7]  ( .D(n3033), .CK(clk), .Q(n4431), 
        .QN(n367) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[6]  ( .D(n3034), .CK(clk), .Q(n4432), 
        .QN(n366) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[8]  ( .D(n3002), .CK(clk), .Q(
        \dp/npc_id_exe_int[8] ), .QN(n4216) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[5]  ( .D(n3035), .CK(clk), .Q(n4433), 
        .QN(n365) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[7]  ( .D(n3003), .CK(clk), .Q(
        \dp/npc_id_exe_int[7] ), .QN(n4210) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[4]  ( .D(n3036), .CK(clk), .Q(n4434), 
        .QN(n364) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[6]  ( .D(n3004), .CK(clk), .Q(
        \dp/npc_id_exe_int[6] ), .QN(n4215) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[3]  ( .D(n3037), .CK(clk), .Q(n4435), 
        .QN(n363) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[5]  ( .D(n3005), .CK(clk), .Q(
        \dp/npc_id_exe_int[5] ), .QN(n4209) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[2]  ( .D(n3038), .CK(clk), .Q(n4412), 
        .QN(n362) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[4]  ( .D(n3006), .CK(clk), .Q(
        \dp/npc_id_exe_int[4] ), .QN(n4214) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[1]  ( .D(n3039), .CK(clk), .Q(n4413), 
        .QN(n361) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[3]  ( .D(n3007), .CK(clk), .Q(
        \dp/npc_id_exe_int[3] ), .QN(n4213) );
  DFF_X1 \dp/ifs/pc/q_reg[0]  ( .D(n2557), .CK(clk), .Q(
        btb_cache_read_address[0]) );
  DFF_X1 \dp/if_id_regs/npc_reg/q_reg[0]  ( .D(n3040), .CK(clk), .Q(n4414), 
        .QN(n360) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[2]  ( .D(n3008), .CK(clk), .Q(
        \dp/npc_id_exe_int[2] ), .QN(btb_cache_rw_address[0]) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[2]  ( .D(n2754), .CK(clk), .Q(
        \dp/op_b_id_ex_int[2] ) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[2]  ( .D(n2619), .CK(clk), .Q(
        dcache_data_out[2]), .QN(n4165) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[2]  ( .D(n2587), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[2] ), .QN(n4441) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[2]  ( .D(n1474), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[2] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[2]  ( .D(n2651), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[2] ), .QN(n4087) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[0]  ( .D(n2653), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[0] ), .QN(n4377) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[0]  ( .D(n2589), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[0] ), .QN(n4440) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[0]  ( .D(n1493), .CK(clk), .Q(
        n4239), .QN(\dp/a_neg_mult_id_exe_int[0] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[31]  ( .D(n2787), .CK(clk), 
        .QN(n681) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[31]  ( .D(n2755), .CK(clk), .Q(
        wp_alu_data_high[31]), .QN(n4539) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[0]  ( .D(n2685), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[0] ) );
  DFF_X1 \dp/id_exe_regs/b10_1_reg/q_reg[1]  ( .D(n2723), .CK(clk), .Q(
        \dp/b10_1_mult_id_exe_int[1] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[1]  ( .D(n2684), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[1] ) );
  DFF_X1 \dp/id_exe_regs/b10_1_reg/q_reg[2]  ( .D(n2722), .CK(clk), .Q(n4231), 
        .QN(n593) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[2]  ( .D(n2683), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[2] ) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[3]  ( .D(n2753), .CK(clk), .Q(
        \dp/op_b_id_ex_int[3] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[3]  ( .D(n2682), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[3] ) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[4]  ( .D(n2752), .CK(clk), .Q(
        \dp/op_b_id_ex_int[4] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[4]  ( .D(n2681), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[4] ) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[5]  ( .D(n2751), .CK(clk), .Q(
        \dp/op_b_id_ex_int[5] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[5]  ( .D(n2680), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[5] ), .QN(n4330) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[6]  ( .D(n2750), .CK(clk), .Q(
        \dp/op_b_id_ex_int[6] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[6]  ( .D(n2679), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[6] ), .QN(n4340) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[7]  ( .D(n2749), .CK(clk), .Q(
        \dp/op_b_id_ex_int[7] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[7]  ( .D(n2678), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[7] ), .QN(n4341) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[8]  ( .D(n2748), .CK(clk), .Q(
        \dp/op_b_id_ex_int[8] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[8]  ( .D(n2677), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[8] ), .QN(n4348) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[9]  ( .D(n2747), .CK(clk), .Q(
        \dp/op_b_id_ex_int[9] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[9]  ( .D(n2676), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[9] ) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[10]  ( .D(n2746), .CK(clk), .Q(
        \dp/op_b_id_ex_int[10] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[10]  ( .D(n2675), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[10] ), .QN(n4347) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[11]  ( .D(n2745), .CK(clk), .Q(
        \dp/op_b_id_ex_int[11] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[11]  ( .D(n2674), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[11] ) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[12]  ( .D(n2744), .CK(clk), .Q(
        \dp/op_b_id_ex_int[12] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[12]  ( .D(n2673), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[12] ), .QN(n4305) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[13]  ( .D(n2743), .CK(clk), .Q(
        \dp/op_b_id_ex_int[13] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[13]  ( .D(n2672), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[13] ), .QN(n4344) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[14]  ( .D(n2742), .CK(clk), .Q(
        \dp/op_b_id_ex_int[14] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[14]  ( .D(n2671), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[14] ), .QN(n4306) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[15]  ( .D(n2741), .CK(clk), .Q(
        \dp/op_b_id_ex_int[15] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[15]  ( .D(n2670), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[15] ), .QN(n4346) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[16]  ( .D(n2740), .CK(clk), .Q(
        \dp/op_b_id_ex_int[16] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[16]  ( .D(n2669), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[16] ), .QN(n4308) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[17]  ( .D(n2739), .CK(clk), .Q(
        \dp/op_b_id_ex_int[17] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[17]  ( .D(n2668), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[17] ), .QN(n4345) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[18]  ( .D(n2738), .CK(clk), .Q(
        \dp/op_b_id_ex_int[18] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[18]  ( .D(n2667), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[18] ), .QN(n4338) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[19]  ( .D(n2737), .CK(clk), .Q(
        \dp/op_b_id_ex_int[19] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[19]  ( .D(n2666), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[19] ), .QN(n4339) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[20]  ( .D(n2736), .CK(clk), .Q(
        \dp/op_b_id_ex_int[20] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[20]  ( .D(n2665), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[20] ), .QN(n4337) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[21]  ( .D(n2735), .CK(clk), .Q(
        \dp/op_b_id_ex_int[21] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[21]  ( .D(n2664), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[21] ), .QN(n4304) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[22]  ( .D(n2734), .CK(clk), .Q(
        \dp/op_b_id_ex_int[22] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[22]  ( .D(n2663), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[22] ), .QN(n4335) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[23]  ( .D(n2733), .CK(clk), .Q(
        \dp/op_b_id_ex_int[23] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[23]  ( .D(n2662), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[23] ), .QN(n4343) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[24]  ( .D(n2732), .CK(clk), .Q(
        \dp/op_b_id_ex_int[24] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[24]  ( .D(n2661), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[24] ), .QN(n4342) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[25]  ( .D(n2731), .CK(clk), .Q(
        \dp/op_b_id_ex_int[25] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[25]  ( .D(n2660), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[25] ), .QN(n4307) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[26]  ( .D(n2730), .CK(clk), .Q(
        \dp/op_b_id_ex_int[26] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[26]  ( .D(n2659), .CK(clk), .QN(n4291) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[27]  ( .D(n2729), .CK(clk), .Q(
        \dp/op_b_id_ex_int[27] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[27]  ( .D(n2658), .CK(clk), .QN(n4295) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[28]  ( .D(n2728), .CK(clk), .Q(
        \dp/op_b_id_ex_int[28] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[28]  ( .D(n2657), .CK(clk), .QN(n4294) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[29]  ( .D(n2727), .CK(clk), .Q(
        \dp/op_b_id_ex_int[29] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[29]  ( .D(n2656), .CK(clk), .QN(n4293) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[30]  ( .D(n2726), .CK(clk), .Q(
        \dp/op_b_id_ex_int[30] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[30]  ( .D(n2655), .CK(clk), .QN(n4292) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[29]  ( .D(n2687), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[29] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[27]  ( .D(n2689), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[27] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[25]  ( .D(n2691), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[25] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[23]  ( .D(n2693), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[23] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[21]  ( .D(n2695), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[21] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[19]  ( .D(n2697), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[19] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[17]  ( .D(n2699), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[17] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[15]  ( .D(n2701), .CK(clk), 
        .Q(n4395) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[13]  ( .D(n2703), .CK(clk), 
        .Q(n4146) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[11]  ( .D(n2705), .CK(clk), 
        .Q(n4392) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[9]  ( .D(n2707), .CK(clk), 
        .Q(n4145) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[7]  ( .D(n2709), .CK(clk), 
        .Q(n4391) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[5]  ( .D(n2711), .CK(clk), 
        .Q(n4141) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[3]  ( .D(n2713), .CK(clk), 
        .Q(n4393) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[1]  ( .D(n2715), .CK(clk), 
        .Q(n5147), .QN(n595) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[31]  ( .D(n2725), .CK(clk), .Q(
        \dp/op_b_id_ex_int[31] ) );
  DFF_X1 \dp/id_exe_regs/b_add_reg/q_reg[31]  ( .D(n2654), .CK(clk), .Q(
        \dp/b_adder_id_exe_int[31] ), .QN(n4582) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[30]  ( .D(n2686), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[30] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[28]  ( .D(n2688), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[28] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[26]  ( .D(n2690), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[26] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[24]  ( .D(n2692), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[24] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[22]  ( .D(n2694), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[22] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[20]  ( .D(n2696), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[20] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[18]  ( .D(n2698), .CK(clk), 
        .Q(\dp/id_exe_regs/b_mult_reg/q[18] ) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[16]  ( .D(n2700), .CK(clk), 
        .Q(n4394) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[14]  ( .D(n2702), .CK(clk), 
        .Q(n4144) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[12]  ( .D(n2704), .CK(clk), 
        .Q(n4390) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[10]  ( .D(n2706), .CK(clk), 
        .Q(n4143) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[8]  ( .D(n2708), .CK(clk), 
        .Q(n4389) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[6]  ( .D(n2710), .CK(clk), 
        .Q(n4142) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[4]  ( .D(n2712), .CK(clk), 
        .Q(n4388) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[2]  ( .D(n2714), .CK(clk), 
        .Q(\dp/b_mult_id_exe_int[2] ), .QN(n5145) );
  DFF_X1 \dp/id_exe_regs/b_mult_reg/curr_data_reg[0]  ( .D(n2716), .CK(clk), 
        .Q(n5146), .QN(n594) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[0]  ( .D(n2882), .CK(clk), .Q(n4482), 
        .QN(n463) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[1]  ( .D(n2881), .CK(clk), .Q(n4255)
         );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[2]  ( .D(n2880), .CK(clk), .Q(n4469), 
        .QN(n465) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[2]  ( .D(n2944), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[2] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[3]  ( .D(n2879), .CK(clk), .Q(n4468), 
        .QN(n466) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[3]  ( .D(n2943), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[3] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[4]  ( .D(n2878), .CK(clk), .Q(n4467), 
        .QN(n467) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[5]  ( .D(n2877), .CK(clk), .Q(n4285)
         );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[6]  ( .D(n2876), .CK(clk), .Q(n4254)
         );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[6]  ( .D(n2940), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[6] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[7]  ( .D(n2875), .CK(clk), .Q(n4253)
         );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[7]  ( .D(n2939), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[7] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[8]  ( .D(n2874), .CK(clk), .Q(n4466), 
        .QN(n471) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[8]  ( .D(n2938), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[8] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[9]  ( .D(n2873), .CK(clk), .Q(n4465), 
        .QN(n472) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[9]  ( .D(n2937), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[9] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[10]  ( .D(n2872), .CK(clk), .Q(n4464), 
        .QN(n473) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[10]  ( .D(n2936), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[10] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[11]  ( .D(n2871), .CK(clk), .Q(n4463), 
        .QN(n474) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[11]  ( .D(n2935), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[11] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[12]  ( .D(n2870), .CK(clk), .Q(n4252)
         );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[12]  ( .D(n2934), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[12] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[13]  ( .D(n2869), .CK(clk), .Q(n4251)
         );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[13]  ( .D(n2933), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[13] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[14]  ( .D(n2868), .CK(clk), .Q(n4250)
         );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[14]  ( .D(n2932), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[14] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[15]  ( .D(n2867), .CK(clk), .Q(n4462), 
        .QN(n478) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[15]  ( .D(n2931), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[15] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[16]  ( .D(n2866), .CK(clk), .Q(n4461), 
        .QN(n479) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[16]  ( .D(n2930), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[16] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[17]  ( .D(n2865), .CK(clk), .Q(n4460), 
        .QN(n480) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[17]  ( .D(n2929), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[17] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[18]  ( .D(n2864), .CK(clk), .Q(n4249)
         );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[19]  ( .D(n2863), .CK(clk), .Q(n4248)
         );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[20]  ( .D(n2862), .CK(clk), .Q(n4247)
         );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[20]  ( .D(n2926), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[20] ), .QN(n4269) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[21]  ( .D(n2861), .CK(clk), .Q(n4246)
         );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[22]  ( .D(n2860), .CK(clk), .Q(n4245)
         );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[23]  ( .D(n2859), .CK(clk), .Q(n4244)
         );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[24]  ( .D(n2858), .CK(clk), .Q(n4243)
         );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[25]  ( .D(n2857), .CK(clk), .Q(n4242)
         );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[26]  ( .D(n2856), .CK(clk), .Q(n4241)
         );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[26]  ( .D(n2920), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[26] ), .QN(n4274) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[27]  ( .D(n2855), .CK(clk), .Q(n4459), 
        .QN(n490) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[28]  ( .D(n2854), .CK(clk), .Q(n4458), 
        .QN(n491) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[29]  ( .D(n2853), .CK(clk), .Q(n4457), 
        .QN(n492) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[29]  ( .D(n2917), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[29] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[30]  ( .D(n2852), .CK(clk), .Q(n4456), 
        .QN(n493) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[30]  ( .D(n2916), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[30] ) );
  DFF_X1 \dp/id_exe_regs/a_add_reg/q_reg[31]  ( .D(n2851), .CK(clk), .Q(n4455), 
        .QN(n494) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[62]  ( .D(n2884), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[62] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[61]  ( .D(n2885), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[61] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[60]  ( .D(n2886), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[60] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[59]  ( .D(n2887), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[59] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[58]  ( .D(n2888), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[58] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[57]  ( .D(n2889), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[57] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[56]  ( .D(n2890), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[56] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[55]  ( .D(n2891), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[55] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[54]  ( .D(n2892), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[54] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[53]  ( .D(n2893), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[53] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[52]  ( .D(n2894), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[52] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[51]  ( .D(n2895), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[51] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[50]  ( .D(n2896), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[50] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[49]  ( .D(n2897), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[49] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[47]  ( .D(n2899), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[47] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[46]  ( .D(n2900), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[46] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[45]  ( .D(n2901), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[45] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[44]  ( .D(n2902), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[44] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[43]  ( .D(n2903), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[43] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[42]  ( .D(n2904), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[42] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[41]  ( .D(n2905), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[41] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[40]  ( .D(n2906), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[40] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[39]  ( .D(n2907), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[39] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[38]  ( .D(n2908), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[38] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[37]  ( .D(n2909), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[37] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[36]  ( .D(n2910), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[36] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[35]  ( .D(n2911), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[35] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[34]  ( .D(n2912), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[34] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[33]  ( .D(n2913), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[33] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[32]  ( .D(n2914), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[32] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[31]  ( .D(n2915), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[31] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[30]  ( .D(n2788), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[62] ), .QN(n7435) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[30]  ( .D(n2756), .CK(clk), .Q(
        wp_alu_data_high[30]), .QN(n4578) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[62]  ( .D(n2820), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[62] ), .QN(n4585) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[29]  ( .D(n2789), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[61] ), .QN(n4179) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[29]  ( .D(n2757), .CK(clk), .Q(
        wp_alu_data_high[29]), .QN(n4577) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[28]  ( .D(n2790), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[60] ), .QN(n7434) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[28]  ( .D(n2758), .CK(clk), .Q(
        wp_alu_data_high[28]), .QN(n4576) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[60]  ( .D(n2822), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[60] ), .QN(n4451) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[27]  ( .D(n2791), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[59] ), .QN(n4204) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[27]  ( .D(n2759), .CK(clk), .Q(
        wp_alu_data_high[27]), .QN(n4575) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[26]  ( .D(n2792), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[58] ), .QN(n4178) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[26]  ( .D(n2760), .CK(clk), .Q(
        wp_alu_data_high[26]), .QN(n4574) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[25]  ( .D(n2793), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[57] ), .QN(n4177) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[25]  ( .D(n2761), .CK(clk), .Q(
        wp_alu_data_high[25]), .QN(n4573) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[57]  ( .D(n2825), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[57] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[24]  ( .D(n2794), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[56] ), .QN(n4187) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[24]  ( .D(n2762), .CK(clk), .Q(
        wp_alu_data_high[24]), .QN(n4572) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[23]  ( .D(n2795), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[55] ), .QN(n4186) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[23]  ( .D(n2763), .CK(clk), .Q(
        wp_alu_data_high[23]), .QN(n4571) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[55]  ( .D(n2827), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[55] ), .QN(n4385) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[22]  ( .D(n2764), .CK(clk), .Q(
        wp_alu_data_high[22]), .QN(n4570) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[54]  ( .D(n2828), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[54] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[21]  ( .D(n2797), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[53] ), .QN(n4176) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[21]  ( .D(n2765), .CK(clk), .Q(
        wp_alu_data_high[21]), .QN(n4569) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[53]  ( .D(n2829), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[53] ), .QN(n4382) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[20]  ( .D(n2798), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[52] ), .QN(n4175) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[20]  ( .D(n2766), .CK(clk), .Q(
        wp_alu_data_high[20]), .QN(n4568) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[19]  ( .D(n2799), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[51] ), .QN(n4194) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[19]  ( .D(n2767), .CK(clk), .Q(
        wp_alu_data_high[19]), .QN(n4567) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[18]  ( .D(n2800), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[50] ), .QN(n7433) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[18]  ( .D(n2768), .CK(clk), .Q(
        wp_alu_data_high[18]), .QN(n4566) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[50]  ( .D(n2832), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[50] ), .QN(n4407) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[17]  ( .D(n2801), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[49] ), .QN(n4193) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[17]  ( .D(n2769), .CK(clk), .Q(
        wp_alu_data_high[17]), .QN(n4565) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[49]  ( .D(n2833), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[49] ), .QN(n4488) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[16]  ( .D(n2802), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[48] ), .QN(n4192) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[16]  ( .D(n2770), .CK(clk), .Q(
        wp_alu_data_high[16]), .QN(n4564) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[48]  ( .D(n2834), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[48] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[15]  ( .D(n2803), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[47] ), .QN(n4191) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[15]  ( .D(n2771), .CK(clk), .Q(
        wp_alu_data_high[15]), .QN(n4563) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[47]  ( .D(n2835), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[47] ), .QN(n4487) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[14]  ( .D(n2804), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[46] ), .QN(n7432) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[14]  ( .D(n2772), .CK(clk), .Q(
        wp_alu_data_high[14]), .QN(n4562) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[46]  ( .D(n2836), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[46] ), .QN(n4486) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[13]  ( .D(n2805), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[45] ), .QN(n4174) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[13]  ( .D(n2773), .CK(clk), .Q(
        wp_alu_data_high[13]), .QN(n4561) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[45]  ( .D(n2837), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[45] ), .QN(n4406) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[12]  ( .D(n2806), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[44] ), .QN(n4173) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[12]  ( .D(n2774), .CK(clk), .Q(
        wp_alu_data_high[12]), .QN(n4560) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[11]  ( .D(n2807), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[43] ), .QN(n4185) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[11]  ( .D(n2775), .CK(clk), .Q(
        wp_alu_data_high[11]), .QN(n4559) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[43]  ( .D(n2839), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[43] ), .QN(n4475) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[10]  ( .D(n2808), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[42] ), .QN(n4184) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[10]  ( .D(n2776), .CK(clk), .Q(
        wp_alu_data_high[10]), .QN(n4558) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[42]  ( .D(n2840), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[42] ), .QN(n4471) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[9]  ( .D(n2809), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[41] ), .QN(n4190) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[9]  ( .D(n2777), .CK(clk), .Q(
        wp_alu_data_high[9]), .QN(n4557) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[41]  ( .D(n2841), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[41] ), .QN(n4504) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[8]  ( .D(n2810), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[40] ), .QN(n7431) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[8]  ( .D(n2778), .CK(clk), .Q(
        wp_alu_data_high[8]), .QN(n4556) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[40]  ( .D(n2842), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[40] ), .QN(n4505) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[7]  ( .D(n2811), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[39] ), .QN(n4189) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[7]  ( .D(n2779), .CK(clk), .Q(
        wp_alu_data_high[7]), .QN(n4555) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[39]  ( .D(n2843), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[39] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[6]  ( .D(n2812), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[38] ), .QN(n4183) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[6]  ( .D(n2780), .CK(clk), .Q(
        wp_alu_data_high[6]), .QN(n4554) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[5]  ( .D(n2813), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[37] ), .QN(n4172) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[5]  ( .D(n2781), .CK(clk), .Q(
        wp_alu_data_high[5]), .QN(n4553) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[4]  ( .D(n2814), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[36] ), .QN(n4171) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[4]  ( .D(n2782), .CK(clk), .Q(
        wp_alu_data_high[4]), .QN(n4552) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[36]  ( .D(n2846), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[36] ), .QN(n4472) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[3]  ( .D(n2815), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[35] ), .QN(n4170) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[3]  ( .D(n2783), .CK(clk), .Q(
        wp_alu_data_high[3]), .QN(n4551) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[35]  ( .D(n2847), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[35] ), .QN(n4453) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[2]  ( .D(n2816), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[34] ), .QN(n7430) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[2]  ( .D(n2784), .CK(clk), .Q(
        wp_alu_data_high[2]), .QN(n4550) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[34]  ( .D(n2848), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[34] ), .QN(n4480) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[1]  ( .D(n2817), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[33] ), .QN(n4188) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[1]  ( .D(n2785), .CK(clk), .Q(
        wp_alu_data_high[1]), .QN(n4549) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[0]  ( .D(n2818), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[32] ), .QN(n4169) );
  DFF_X1 \dp/mem_wb_regs/alu_high_reg/q_reg[0]  ( .D(n2786), .CK(clk), .Q(
        wp_alu_data_high[0]), .QN(n4548) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[32]  ( .D(n2850), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[32] ), .QN(n4403) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[1]  ( .D(n1475), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[1] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[1]  ( .D(n2652), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[1] ), .QN(n4072) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[1]  ( .D(n2588), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[1] ), .QN(n4439) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[1]  ( .D(n2620), .CK(clk), .Q(
        dcache_data_out[1]), .QN(n4163) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[3]  ( .D(n1473), .CK(clk), .Q(
        n4227), .QN(\dp/a_neg_mult_id_exe_int[3] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[3]  ( .D(n2650), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[3] ), .QN(n4080) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[3]  ( .D(n2586), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[3] ), .QN(n4438) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[3]  ( .D(n2618), .CK(clk), .Q(
        dcache_data_out[3]), .QN(n4162) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[4]  ( .D(n1472), .CK(clk), .Q(
        n4105), .QN(\dp/a_neg_mult_id_exe_int[4] ) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[4]  ( .D(n2585), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[4] ), .QN(n4437) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[4]  ( .D(n2617), .CK(clk), .Q(
        dcache_data_out[4]), .QN(n4161) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[5]  ( .D(n2648), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[5] ), .QN(n6459) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[5]  ( .D(n2584), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[5] ), .QN(n4516) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[5]  ( .D(n2616), .CK(clk), .Q(
        dcache_data_out[5]), .QN(n4160) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[6]  ( .D(n1470), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[6] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[6]  ( .D(n2647), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[6] ), .QN(n6456) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[6]  ( .D(n2583), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[6] ), .QN(n4515) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[6]  ( .D(n2615), .CK(clk), .Q(
        dcache_data_out[6]), .QN(n4159) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[7]  ( .D(n1469), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[7] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[7]  ( .D(n2646), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[7] ), .QN(n6453) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[7]  ( .D(n2582), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[7] ), .QN(n4514) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[7]  ( .D(n2614), .CK(clk), .Q(
        dcache_data_out[7]), .QN(n4158) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[8]  ( .D(n1468), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[8] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[8]  ( .D(n2645), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[8] ), .QN(n4063) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[8]  ( .D(n2581), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[8] ), .QN(n4513) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[8]  ( .D(n2613), .CK(clk), .Q(
        dcache_data_out[8]), .QN(n4157) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[9]  ( .D(n1467), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[9] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[9]  ( .D(n2644), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[9] ), .QN(n4082) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[9]  ( .D(n2580), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[9] ), .QN(n4512) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[9]  ( .D(n2612), .CK(clk), .Q(
        dcache_data_out[9]), .QN(n4156) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[10]  ( .D(n1466), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[10] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[10]  ( .D(n2643), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[10] ), .QN(n4074) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[10]  ( .D(n2579), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[10] ), .QN(n4511) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[10]  ( .D(n2611), .CK(clk), .Q(
        dcache_data_out[10]), .QN(n4155) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[11]  ( .D(n1465), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[11] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[11]  ( .D(n2642), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[11] ), .QN(n4073) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[11]  ( .D(n2578), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[11] ), .QN(n4510) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[11]  ( .D(n2610), .CK(clk), .Q(
        dcache_data_out[11]), .QN(n4154) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[12]  ( .D(n1464), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[12] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[12]  ( .D(n2641), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[12] ), .QN(n4088) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[12]  ( .D(n2577), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[12] ), .QN(n4509) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[12]  ( .D(n2609), .CK(clk), .Q(
        dcache_data_out[12]), .QN(n4153) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[13]  ( .D(n1463), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[13] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[13]  ( .D(n2640), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[13] ), .QN(n4079) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[13]  ( .D(n2576), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[13] ), .QN(n4508) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[13]  ( .D(n2608), .CK(clk), .Q(
        dcache_data_out[13]), .QN(n4152) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[14]  ( .D(n1462), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[14] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[14]  ( .D(n2639), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[14] ), .QN(n4066) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[14]  ( .D(n2575), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[14] ), .QN(n4507) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[14]  ( .D(n2607), .CK(clk), .Q(
        dcache_data_out[14]), .QN(n4151) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[15]  ( .D(n2638), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[15] ), .QN(n4081) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[15]  ( .D(n2574), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[15] ), .QN(n4506) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[15]  ( .D(n2606), .CK(clk), .Q(
        dcache_data_out[15]), .QN(n4150) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[16]  ( .D(n2637), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[16] ), .QN(n4089) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[16]  ( .D(n2573), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[16] ), .QN(n4587) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[16]  ( .D(n2605), .CK(clk), .Q(
        dcache_data_out[16]), .QN(n4196) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[17]  ( .D(n2636), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[17] ), .QN(n4095) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[17]  ( .D(n2572), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[17] ), .QN(n4588) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[17]  ( .D(n2604), .CK(clk), .Q(
        dcache_data_out[17]), .QN(n4197) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[18]  ( .D(n2635), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[18] ), .QN(n4085) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[18]  ( .D(n2571), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[18] ), .QN(n4589) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[18]  ( .D(n2603), .CK(clk), .Q(
        dcache_data_out[18]), .QN(n4198) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[19]  ( .D(n2634), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[19] ), .QN(n4075) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[19]  ( .D(n2570), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[19] ), .QN(n4590) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[19]  ( .D(n2602), .CK(clk), .Q(
        dcache_data_out[19]), .QN(n4199) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[20]  ( .D(n2633), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[20] ), .QN(n4076) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[20]  ( .D(n2569), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[20] ), .QN(n4591) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[20]  ( .D(n2601), .CK(clk), .Q(
        dcache_data_out[20]), .QN(n4200) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[21]  ( .D(n2632), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[21] ), .QN(n4086) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[21]  ( .D(n2568), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[21] ), .QN(n4592) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[21]  ( .D(n2600), .CK(clk), .Q(
        dcache_data_out[21]), .QN(n4201) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[22]  ( .D(n1454), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[22] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[22]  ( .D(n2631), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[22] ), .QN(n4077) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[22]  ( .D(n2567), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[22] ), .QN(n4593) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[22]  ( .D(n2599), .CK(clk), .Q(
        dcache_data_out[22]), .QN(n4202) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[23]  ( .D(n1453), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[23] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[23]  ( .D(n2630), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[23] ), .QN(n4078) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[23]  ( .D(n2566), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[23] ), .QN(n4594) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[23]  ( .D(n2598), .CK(clk), .Q(
        dcache_data_out[23]), .QN(n4203) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[24]  ( .D(n1452), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[24] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[24]  ( .D(n2629), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[24] ), .QN(n4084) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[24]  ( .D(n2565), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[24] ), .QN(n4112) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[24]  ( .D(n2597), .CK(clk), .Q(
        dcache_data_out[24]), .QN(n4530) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[25]  ( .D(n1451), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[25] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[25]  ( .D(n2628), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[25] ), .QN(n4062) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[25]  ( .D(n2564), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[25] ), .QN(n4090) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[25]  ( .D(n2596), .CK(clk), .Q(
        dcache_data_out[25]), .QN(n4531) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[26]  ( .D(n1450), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[26] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[26]  ( .D(n2627), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[26] ), .QN(n4065) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[26]  ( .D(n2563), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[26] ), .QN(n4091) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[26]  ( .D(n2595), .CK(clk), .Q(
        dcache_data_out[26]), .QN(n4532) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[27]  ( .D(n1449), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[27] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[27]  ( .D(n2626), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[27] ), .QN(n4064) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[27]  ( .D(n2562), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[27] ), .QN(n4092) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[27]  ( .D(n2594), .CK(clk), .Q(
        dcache_data_out[27]), .QN(n4533) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[28]  ( .D(n1448), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[28] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[28]  ( .D(n2625), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[28] ), .QN(n4067) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[28]  ( .D(n2561), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[28] ), .QN(n4093) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[28]  ( .D(n2593), .CK(clk), .Q(
        dcache_data_out[28]), .QN(n4534) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[29]  ( .D(n1447), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[29] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[29]  ( .D(n2624), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[29] ), .QN(n4068) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[29]  ( .D(n2560), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[29] ), .QN(n4094) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[29]  ( .D(n2592), .CK(clk), .Q(
        dcache_data_out[29]), .QN(n4535) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[30]  ( .D(n1446), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[30] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[30]  ( .D(n2623), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[30] ), .QN(n4109) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[30]  ( .D(n2559), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[30] ), .QN(n7496) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[30]  ( .D(n2591), .CK(clk), .Q(
        dcache_data_out[30]), .QN(n4401) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[31]  ( .D(n1444), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[31] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[31]  ( .D(n2622), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[31] ), .QN(n4096) );
  DFF_X1 \dp/mem_wb_regs/alu_low_reg/q_reg[31]  ( .D(n2558), .CK(clk), .Q(
        \dp/alu_out_low_mem_wb_int[31] ), .QN(n4436) );
  DFF_X1 \dp/ifs/pc/q_reg[27]  ( .D(n2530), .CK(clk), .Q(
        btb_cache_read_address[27]) );
  DFF_X1 \dp/ifs/pc/q_reg[26]  ( .D(n2531), .CK(clk), .Q(
        btb_cache_read_address[26]), .QN(n4598) );
  DFF_X1 \dp/ifs/pc/q_reg[24]  ( .D(n2533), .CK(clk), .Q(
        btb_cache_read_address[24]), .QN(n4597) );
  DFF_X1 \dp/ifs/pc/q_reg[23]  ( .D(n2534), .CK(clk), .Q(
        btb_cache_read_address[23]), .QN(n4596) );
  DFF_X1 \dp/ifs/pc/q_reg[22]  ( .D(n2535), .CK(clk), .Q(
        btb_cache_read_address[22]) );
  DFF_X1 \dp/ifs/pc/q_reg[21]  ( .D(n2536), .CK(clk), .Q(
        btb_cache_read_address[21]) );
  DFF_X1 \dp/ifs/pc/q_reg[20]  ( .D(n2537), .CK(clk), .Q(
        btb_cache_read_address[20]) );
  DFF_X1 \dp/ifs/pc/q_reg[19]  ( .D(n2538), .CK(clk), .Q(
        btb_cache_read_address[19]) );
  DFF_X1 \dp/ifs/pc/q_reg[18]  ( .D(n2539), .CK(clk), .Q(
        btb_cache_read_address[18]) );
  DFF_X1 \dp/ifs/pc/q_reg[17]  ( .D(n2540), .CK(clk), .Q(
        btb_cache_read_address[17]) );
  DFF_X1 \dp/ifs/pc/q_reg[16]  ( .D(n2541), .CK(clk), .Q(
        btb_cache_read_address[16]) );
  DFF_X1 \dp/ifs/pc/q_reg[15]  ( .D(n2542), .CK(clk), .Q(
        btb_cache_read_address[15]) );
  DFF_X1 \dp/ifs/pc/q_reg[14]  ( .D(n2543), .CK(clk), .Q(
        btb_cache_read_address[14]) );
  DFF_X1 \dp/ifs/pc/q_reg[13]  ( .D(n2544), .CK(clk), .Q(
        btb_cache_read_address[13]) );
  DFF_X1 \dp/ifs/pc/q_reg[12]  ( .D(n2545), .CK(clk), .Q(
        btb_cache_read_address[12]) );
  DFF_X1 \dp/ifs/pc/q_reg[11]  ( .D(n2546), .CK(clk), .Q(
        btb_cache_read_address[11]) );
  DFF_X1 \dp/ifs/pc/q_reg[10]  ( .D(n2547), .CK(clk), .Q(
        btb_cache_read_address[10]) );
  DFF_X1 \dp/ifs/pc/q_reg[9]  ( .D(n2548), .CK(clk), .Q(
        btb_cache_read_address[9]) );
  DFF_X1 \dp/ifs/pc/q_reg[8]  ( .D(n2549), .CK(clk), .Q(
        btb_cache_read_address[8]) );
  DFF_X1 \dp/ifs/pc/q_reg[7]  ( .D(n2550), .CK(clk), .Q(
        btb_cache_read_address[7]) );
  DFF_X1 \dp/ifs/pc/q_reg[6]  ( .D(n2551), .CK(clk), .Q(
        btb_cache_read_address[6]) );
  DFF_X1 \dp/ifs/pc/q_reg[5]  ( .D(n2552), .CK(clk), .Q(
        btb_cache_read_address[5]) );
  DFF_X1 \dp/ifs/pc/q_reg[4]  ( .D(n2553), .CK(clk), .Q(
        btb_cache_read_address[4]) );
  DFF_X1 \dp/ifs/pc/q_reg[3]  ( .D(n2554), .CK(clk), .Q(
        btb_cache_read_address[3]) );
  DFF_X1 \dp/ifs/pc/q_reg[2]  ( .D(n2555), .CK(clk), .Q(
        btb_cache_read_address[2]), .QN(n3868) );
  DFF_X1 \dp/ifs/pc/q_reg[1]  ( .D(n2556), .CK(clk), .Q(
        btb_cache_read_address[1]) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[31]  ( .D(n2590), .CK(clk), .Q(
        dcache_data_out[31]), .QN(n4149) );
  DFF_X1 \dp/ex_mem_regs/b_reg/q_reg[0]  ( .D(n2621), .CK(clk), .Q(
        dcache_data_out[0]), .QN(n4164) );
  DFF_X1 \dp/ifs/pc/q_reg[29]  ( .D(n3041), .CK(clk), .Q(
        btb_cache_read_address[29]), .QN(n3966) );
  DFF_X1 \ctrl_u/curr_id_reg[25]  ( .D(\ctrl_u/n335 ), .CK(clk), .Q(n4478), 
        .QN(\ctrl_u/curr_id[25] ) );
  DFF_X1 \ctrl_u/curr_id_reg[23]  ( .D(\ctrl_u/n535 ), .CK(clk), .QN(n4492) );
  DFF_X1 \ctrl_u/curr_mul_id_reg  ( .D(\ctrl_u/n69 ), .CK(clk), .Q(n4318), 
        .QN(\ctrl_u/n83 ) );
  DFF_X1 \ctrl_u/curr_id_reg[17]  ( .D(\ctrl_u/n541 ), .CK(clk), .Q(
        \ctrl_u/curr_id[17] ), .QN(n4484) );
  DFF_X1 \ctrl_u/curr_id_reg[18]  ( .D(\ctrl_u/n540 ), .CK(clk), .Q(
        \ctrl_u/curr_id[18] ), .QN(\ctrl_u/n70 ) );
  DFF_X1 \ctrl_u/curr_id_reg[6]  ( .D(\ctrl_u/n402 ), .CK(clk), .QN(
        \ctrl_u/curr_id[6] ) );
  DFF_X1 \ctrl_u/curr_id_reg[2]  ( .D(\ctrl_u/n552 ), .CK(clk), .Q(
        \ctrl_u/curr_id[2] ), .QN(\ctrl_u/n74 ) );
  DFF_X1 \ctrl_u/curr_id_reg[3]  ( .D(\ctrl_u/n551 ), .CK(clk), .Q(
        \ctrl_u/curr_id[3] ), .QN(\ctrl_u/n73 ) );
  DFF_X1 \ctrl_u/curr_id_reg[4]  ( .D(\ctrl_u/n550 ), .CK(clk), .Q(
        \ctrl_u/curr_id[4] ), .QN(\ctrl_u/n72 ) );
  DFF_X1 \ctrl_u/curr_id_reg[15]  ( .D(\ctrl_u/n543 ), .CK(clk), .QN(n4454) );
  DFF_X1 \ctrl_u/curr_id_reg[45]  ( .D(\ctrl_u/n518 ), .CK(clk), .QN(
        \ctrl_u/n66 ) );
  DFF_X1 \ctrl_u/curr_id_reg[51]  ( .D(\ctrl_u/n512 ), .CK(clk), .Q(n4481), 
        .QN(\ctrl_u/n62 ) );
  DFF_X1 \ctrl_u/curr_id_reg[50]  ( .D(\ctrl_u/n513 ), .CK(clk), .QN(
        \ctrl_u/n63 ) );
  DFF_X1 \ctrl_u/curr_id_reg[46]  ( .D(\ctrl_u/n517 ), .CK(clk), .QN(
        \ctrl_u/n65 ) );
  DFF_X1 \ctrl_u/curr_id_reg[44]  ( .D(\ctrl_u/n519 ), .CK(clk), .QN(
        \ctrl_u/n67 ) );
  DFF_X1 \ctrl_u/curr_id_reg[43]  ( .D(\ctrl_u/n520 ), .CK(clk), .QN(
        \ctrl_u/n68 ) );
  DFF_X1 \ctrl_u/curr_id_reg[62]  ( .D(\ctrl_u/n554 ), .CK(clk), .QN(n4396) );
  DFF_X1 \ctrl_u/curr_id_reg[1]  ( .D(\ctrl_u/n412 ), .CK(clk), .QN(
        \ctrl_u/curr_id[1] ) );
  DFF_X1 \ctrl_u/curr_id_reg[5]  ( .D(\ctrl_u/n406 ), .CK(clk), .QN(
        \ctrl_u/curr_id[5] ) );
  DFF_X1 \ctrl_u/curr_id_reg[8]  ( .D(\ctrl_u/n548 ), .CK(clk), .Q(
        \ctrl_u/curr_id[8] ), .QN(n4543) );
  DFF_X1 \ctrl_u/curr_id_reg[9]  ( .D(\ctrl_u/n547 ), .CK(clk), .Q(
        \ctrl_u/curr_id[9] ), .QN(n4542) );
  DFF_X1 \ctrl_u/curr_id_reg[10]  ( .D(\ctrl_u/n546 ), .CK(clk), .Q(
        \ctrl_u/curr_id[10] ), .QN(n4541) );
  DFF_X1 \ctrl_u/curr_id_reg[11]  ( .D(\ctrl_u/n545 ), .CK(clk), .Q(
        \ctrl_u/curr_id[11] ), .QN(n4540) );
  DFF_X1 \ctrl_u/curr_id_reg[13]  ( .D(\ctrl_u/n386 ), .CK(clk), .QN(
        \ctrl_u/curr_id[13] ) );
  DFF_X1 \ctrl_u/curr_id_reg[14]  ( .D(\ctrl_u/n384 ), .CK(clk), .QN(
        \ctrl_u/curr_id[14] ) );
  DFF_X1 \ctrl_u/curr_id_reg[19]  ( .D(\ctrl_u/n539 ), .CK(clk), .Q(
        \ctrl_u/curr_id[19] ), .QN(n4546) );
  DFF_X1 \ctrl_u/curr_id_reg[20]  ( .D(\ctrl_u/n538 ), .CK(clk), .Q(
        \ctrl_u/curr_id[20] ), .QN(n4545) );
  DFF_X1 \ctrl_u/curr_id_reg[21]  ( .D(\ctrl_u/n537 ), .CK(clk), .Q(
        \ctrl_u/curr_id[21] ), .QN(n4544) );
  DFF_X1 \ctrl_u/curr_id_reg[27]  ( .D(\ctrl_u/n532 ), .CK(clk), .Q(
        \ctrl_u/curr_id[27] ), .QN(n4581) );
  DFF_X1 \ctrl_u/curr_id_reg[31]  ( .D(\ctrl_u/n305 ), .CK(clk), .QN(
        \ctrl_u/curr_id[31] ) );
  DFF_X1 \ctrl_u/curr_id_reg[32]  ( .D(\ctrl_u/n303 ), .CK(clk), .QN(
        \ctrl_u/curr_id[32] ) );
  DFF_X1 \ctrl_u/curr_id_reg[33]  ( .D(\ctrl_u/n301 ), .CK(clk), .QN(
        \ctrl_u/curr_id[33] ) );
  DFF_X1 \ctrl_u/curr_id_reg[36]  ( .D(\ctrl_u/n526 ), .CK(clk), .Q(
        \ctrl_u/curr_id[36] ), .QN(n4600) );
  DFF_X1 \ctrl_u/curr_id_reg[38]  ( .D(\ctrl_u/n524 ), .CK(clk), .Q(
        \ctrl_u/curr_id[38] ), .QN(n4601) );
  DFF_X1 \ctrl_u/curr_id_reg[40]  ( .D(\ctrl_u/n245 ), .CK(clk), .QN(
        \ctrl_u/curr_id[40] ) );
  DFF_X1 \ctrl_u/curr_id_reg[41]  ( .D(\ctrl_u/n522 ), .CK(clk), .Q(
        \ctrl_u/curr_id[41] ), .QN(n4580) );
  DFF_X1 \ctrl_u/curr_id_reg[52]  ( .D(\ctrl_u/n511 ), .CK(clk), .Q(
        data_tbs_selector_id), .QN(n4584) );
  DFF_X1 \ctrl_u/curr_id_reg[56]  ( .D(\ctrl_u/n508 ), .CK(clk), .Q(
        is_signed_id), .QN(n4502) );
  DFF_X1 \ctrl_u/curr_id_reg[57]  ( .D(\ctrl_u/n181 ), .CK(clk), .QN(
        rp2_out_sel_id[0]) );
  DFF_X1 \ctrl_u/curr_id_reg[58]  ( .D(\ctrl_u/n179 ), .CK(clk), .QN(
        rp2_out_sel_id[1]) );
  DFF_X1 \ctrl_u/curr_id_reg[61]  ( .D(\ctrl_u/n505 ), .CK(clk), .Q(j_instr_id), .QN(n4579) );
  DFF_X1 \ctrl_u/curr_id_reg[29]  ( .D(\ctrl_u/n530 ), .CK(clk), .Q(
        \ctrl_u/curr_id[29] ), .QN(\ctrl_u/n59 ) );
  DFF_X1 \ctrl_u/curr_id_reg[26]  ( .D(\ctrl_u/n533 ), .CK(clk), .Q(
        \ctrl_u/curr_id[26] ), .QN(\ctrl_u/n61 ) );
  DFF_X1 \ctrl_u/curr_id_reg[49]  ( .D(\ctrl_u/n514 ), .CK(clk), .Q(n4485), 
        .QN(\ctrl_u/n64 ) );
  DFF_X1 \ctrl_u/curr_id_reg[34]  ( .D(\ctrl_u/n528 ), .CK(clk), .Q(
        \ctrl_u/curr_id[34] ), .QN(n4521) );
  DFF_X1 \ctrl_u/curr_id_reg[24]  ( .D(\ctrl_u/n534 ), .CK(clk), .QN(n4491) );
  DFF_X1 \ctrl_u/curr_id_reg[35]  ( .D(\ctrl_u/n527 ), .CK(clk), .Q(
        \ctrl_u/curr_id[35] ), .QN(n4522) );
  DFF_X1 \ctrl_u/curr_id_reg[7]  ( .D(\ctrl_u/n549 ), .CK(clk), .Q(
        \ctrl_u/curr_id[7] ), .QN(n4602) );
  DFF_X1 \ctrl_u/curr_id_reg[16]  ( .D(\ctrl_u/n542 ), .CK(clk), .Q(
        \ctrl_u/curr_id[16] ), .QN(n4586) );
  DFF_X1 \ctrl_u/curr_id_reg[42]  ( .D(\ctrl_u/n521 ), .CK(clk), .QN(n4547) );
  DFF_X1 \ctrl_u/curr_ak_exe_reg  ( .D(\ctrl_u/n169 ), .CK(clk), .QN(
        \ctrl_u/curr_ak_exe ) );
  DFF_X1 \ctrl_u/curr_ak_id_reg  ( .D(\ctrl_u/n170 ), .CK(clk), .QN(
        \ctrl_u/curr_ak_id ) );
  DFF_X1 \ctrl_u/curr_pt_exe_reg  ( .D(\ctrl_u/n166 ), .CK(clk), .QN(
        \ctrl_u/curr_pt_exe ) );
  DFF_X1 \ctrl_u/curr_pt_id_reg  ( .D(\ctrl_u/n167 ), .CK(clk), .QN(
        \ctrl_u/curr_pt_id ) );
  DFF_X1 \ctrl_u/curr_exe_reg[29]  ( .D(\ctrl_u/n432 ), .CK(clk), .Q(
        op_type_exe[1]), .QN(\ctrl_u/op_type_exe[1] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[22]  ( .D(\ctrl_u/n439 ), .CK(clk), .QN(
        alu_comp_sel[1]) );
  DFF_X1 \ctrl_u/curr_exe_reg[18]  ( .D(\ctrl_u/n443 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[18] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[6]  ( .D(\ctrl_u/n455 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[6] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[4]  ( .D(\ctrl_u/n457 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[4] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[3]  ( .D(\ctrl_u/n458 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[3] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[2]  ( .D(\ctrl_u/n459 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[2] ) );
  DFF_X1 \ctrl_u/curr_it_reg[2]  ( .D(\ctrl_u/n501 ), .CK(clk), .Q(it_exe[2]), 
        .QN(n5161) );
  DFF_X1 \ctrl_u/curr_it_reg[0]  ( .D(\ctrl_u/n503 ), .CK(clk), .Q(n5159), 
        .QN(n5165) );
  DFF_X1 \ctrl_u/curr_it_reg[3]  ( .D(\ctrl_u/n504 ), .CK(clk), .Q(it_exe[3]), 
        .QN(n5148) );
  DFF_X1 \ctrl_u/curr_it_reg[1]  ( .D(\ctrl_u/n502 ), .CK(clk), .Q(it_exe[1]), 
        .QN(n5163) );
  DFF_X1 \ctrl_u/curr_es_reg[1]  ( .D(\ctrl_u/n558 ), .CK(clk), .Q(n5157), 
        .QN(\ctrl_u/n94 ) );
  DFF_X1 \ctrl_u/curr_exe_reg[0]  ( .D(\ctrl_u/n461 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[0] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[1]  ( .D(\ctrl_u/n460 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[1] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[5]  ( .D(\ctrl_u/n456 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[5] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[9]  ( .D(\ctrl_u/n452 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[9] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[11]  ( .D(\ctrl_u/n450 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[11] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[12]  ( .D(\ctrl_u/n449 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[12] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[13]  ( .D(\ctrl_u/n448 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[13] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[14]  ( .D(\ctrl_u/n447 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[14] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[16]  ( .D(\ctrl_u/n445 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[16] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[19]  ( .D(\ctrl_u/n442 ), .CK(clk), .QN(
        \ctrl_u/curr_exe[19] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[31]  ( .D(\ctrl_u/n430 ), .CK(clk), .QN(
        log_type_exe[1]) );
  DFF_X1 \ctrl_u/curr_exe_reg[32]  ( .D(\ctrl_u/n429 ), .CK(clk), .QN(
        log_type_exe[2]) );
  DFF_X1 \ctrl_u/curr_exe_reg[33]  ( .D(\ctrl_u/n428 ), .CK(clk), .QN(
        log_type_exe[3]) );
  DFF_X1 \ctrl_u/curr_exe_reg[36]  ( .D(\ctrl_u/n425 ), .CK(clk), .QN(
        shift_type_exe[2]) );
  DFF_X1 \ctrl_u/curr_exe_reg[40]  ( .D(\ctrl_u/n421 ), .CK(clk), .QN(
        \ctrl_u/curr_exe_40 ) );
  DFF_X1 \ctrl_u/curr_exe_reg[41]  ( .D(\ctrl_u/n420 ), .CK(clk), .QN(
        \ctrl_u/curr_exe_41 ) );
  DFF_X1 \ctrl_u/curr_ms_reg  ( .D(\ctrl_u/n555 ), .CK(clk), .Q(
        \ctrl_u/curr_ms ), .QN(n4127) );
  DFF_X1 \ctrl_u/curr_mem_reg[14]  ( .D(\ctrl_u/n465 ), .CK(clk), .QN(
        cpu_is_reading) );
  DFF_X1 \ctrl_u/curr_mem_reg[13]  ( .D(\ctrl_u/n467 ), .CK(clk), .Q(n4303), 
        .QN(wr_mem) );
  DFF_X1 \ctrl_u/curr_mem_reg[12]  ( .D(\ctrl_u/n468 ), .CK(clk), .QN(
        \ctrl_u/curr_mem_12 ) );
  DFF_X1 \ctrl_u/curr_mem_reg[11]  ( .D(\ctrl_u/n469 ), .CK(clk), .QN(
        \ctrl_u/curr_mem_11 ) );
  DFF_X1 \ctrl_u/curr_mem_reg[10]  ( .D(\ctrl_u/n470 ), .CK(clk), .Q(n4166), 
        .QN(ld_sign_mem) );
  DFF_X1 \ctrl_u/curr_mem_reg[9]  ( .D(\ctrl_u/n471 ), .CK(clk), .Q(n4386), 
        .QN(ld_type_mem[1]) );
  DFF_X1 \ctrl_u/curr_mem_reg[8]  ( .D(\ctrl_u/n472 ), .CK(clk), .Q(n4470), 
        .QN(ld_type_mem[0]) );
  DFF_X1 \ctrl_u/curr_mem_reg[7]  ( .D(\ctrl_u/n473 ), .CK(clk), .Q(n4479), 
        .QN(alu_data_tbs_selector) );
  DFF_X1 \ctrl_u/curr_mem_reg[6]  ( .D(\ctrl_u/n474 ), .CK(clk), .QN(
        \ctrl_u/curr_mem[6] ) );
  DFF_X1 \ctrl_u/curr_mem_reg[5]  ( .D(\ctrl_u/n475 ), .CK(clk), .QN(
        \ctrl_u/curr_mem[5] ) );
  DFF_X1 \ctrl_u/curr_mem_reg[4]  ( .D(\ctrl_u/n476 ), .CK(clk), .QN(
        \ctrl_u/curr_mem[4] ) );
  DFF_X1 \ctrl_u/curr_mem_reg[2]  ( .D(\ctrl_u/n478 ), .CK(clk), .QN(
        \ctrl_u/curr_mem[2] ) );
  DFF_X1 \ctrl_u/curr_mem_reg[1]  ( .D(\ctrl_u/n479 ), .CK(clk), .QN(
        \ctrl_u/curr_mem[1] ) );
  DFF_X1 \ctrl_u/curr_mem_reg[0]  ( .D(\ctrl_u/n480 ), .CK(clk), .QN(
        \ctrl_u/curr_mem[0] ) );
  DFF_X1 \ctrl_u/curr_wb_reg[3]  ( .D(\ctrl_u/n481 ), .CK(clk), .QN(
        \ctrl_u/curr_wb[3] ) );
  DFF_X1 \ctrl_u/curr_wb_reg[2]  ( .D(\ctrl_u/n483 ), .CK(clk), .QN(wp_en) );
  DFF_X1 \ctrl_u/curr_wb_reg[0]  ( .D(\ctrl_u/n486 ), .CK(clk), .QN(hilo_wr_en) );
  DFF_X1 \ctrl_u/curr_es_reg[0]  ( .D(\ctrl_u/n557 ), .CK(clk), .Q(n5160), 
        .QN(\ctrl_u/n95 ) );
  DFF_X1 \ctrl_u/curr_mul_end_wb_reg  ( .D(\ctrl_u/n559 ), .CK(clk), .Q(
        \ctrl_u/curr_mul_end_wb ), .QN(n4595) );
  FA_X1 \intadd_2/U23  ( .A(\intadd_2/A[6] ), .B(n4217), .CI(\intadd_2/n23 ), 
        .CO(\intadd_2/n22 ), .S(\intadd_2/SUM[6] ) );
  FA_X1 \intadd_2/U22  ( .A(n4121), .B(n4233), .CI(\intadd_2/n22 ), .CO(
        \intadd_2/n21 ), .S(\intadd_2/SUM[7] ) );
  FA_X1 \intadd_2/U21  ( .A(\intadd_2/A[8] ), .B(n4218), .CI(\intadd_2/n21 ), 
        .CO(\intadd_2/n20 ), .S(\intadd_2/SUM[8] ) );
  FA_X1 \intadd_2/U20  ( .A(n4120), .B(n4234), .CI(\intadd_2/n20 ), .CO(
        \intadd_2/n19 ), .S(\intadd_2/SUM[9] ) );
  FA_X1 \intadd_2/U19  ( .A(n4119), .B(n4226), .CI(\intadd_2/n19 ), .CO(
        \intadd_2/n18 ), .S(\intadd_2/SUM[10] ) );
  FA_X1 \intadd_2/U18  ( .A(n4118), .B(n4235), .CI(\intadd_2/n18 ), .CO(
        \intadd_2/n17 ), .S(\intadd_2/SUM[11] ) );
  FA_X1 \intadd_2/U13  ( .A(n4258), .B(n4110), .CI(\intadd_2/n13 ), .CO(
        \intadd_2/n12 ), .S(\intadd_2/SUM[16] ) );
  FA_X1 \intadd_2/U12  ( .A(n4259), .B(n4114), .CI(\intadd_2/n12 ), .CO(
        \intadd_2/n11 ), .S(\intadd_2/SUM[17] ) );
  FA_X1 \intadd_2/U6  ( .A(n4397), .B(n4147), .CI(\intadd_2/n6 ), .CO(
        \intadd_2/n5 ), .S(\intadd_2/SUM[23] ) );
  FA_X1 \intadd_2/U5  ( .A(n4398), .B(n4520), .CI(\intadd_2/n5 ), .CO(
        \intadd_2/n4 ), .S(\intadd_2/SUM[24] ) );
  FA_X1 \intadd_2/U4  ( .A(n4399), .B(n4148), .CI(\intadd_2/n4 ), .CO(
        \intadd_2/n3 ), .S(\intadd_2/SUM[25] ) );
  FA_X1 \intadd_2/U3  ( .A(n4400), .B(n4536), .CI(\intadd_2/n3 ), .CO(
        \intadd_2/n2 ), .S(\intadd_2/SUM[26] ) );
  DFF_X2 \ctrl_u/curr_mul_in_prog_reg  ( .D(\ctrl_u/n556 ), .CK(clk), .Q(
        \ctrl_u/curr_mul_in_prog ), .QN(n4238) );
  DFF_X2 \ctrl_u/curr_exe_reg[38]  ( .D(\ctrl_u/n423 ), .CK(clk), .Q(n4225), 
        .QN(sub_add_exe) );
  TBUF_X1 \ctrl_u/en_npc_id_tri2  ( .A(1'b0), .EN(n3933), .Z(en_npc_id) );
  TBUF_X1 \ctrl_u/en_rd_id_tri2  ( .A(1'b0), .EN(n3933), .Z(en_rd_id) );
  TBUF_X1 \ctrl_u/en_shift_id_tri2  ( .A(1'b0), .EN(n3933), .Z(en_shift_id) );
  TBUF_X1 \ctrl_u/en_imm_id_tri2  ( .A(1'b0), .EN(n3933), .Z(en_imm_id) );
  TBUF_X1 \ctrl_u/en_shift_reg_id_tri2  ( .A(n7274), .EN(n3933), .Z(
        en_shift_reg_id) );
  TBUF_X1 \ctrl_u/en_b_id_tri2  ( .A(1'b0), .EN(n3933), .Z(en_b_id) );
  TBUF_X1 \ctrl_u/en_mul_id_tri2  ( .A(1'b0), .EN(n3933), .Z(en_mul_id) );
  TBUF_X1 \ctrl_u/en_add_id_tri2  ( .A(1'b0), .EN(n3933), .Z(en_add_id) );
  TBUF_X1 \ctrl_u/shift_reg_id_tri2  ( .A(n7274), .EN(n3933), .Z(shift_reg_id)
         );
  TBUF_X1 \mc/cache_update_type_tri[1]  ( .A(1'b0), .EN(n3910), .Z(
        dcache_update_type[1]) );
  TBUF_X1 \mc/cache_update_type_tri[0]  ( .A(1'b0), .EN(n3910), .Z(
        dcache_update_type[0]) );
  TBUF_X1 \mc/cache_update_tri  ( .A(1'b1), .EN(n3910), .Z(dcache_update) );
  TBUF_X1 \ctrl_u/dcache_update_tri  ( .A(wr_mem), .EN(\ctrl_u/curr_ms ), .Z(
        dcache_update) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[59]  ( .D(n2823), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[59] ), .QN(n4537) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[22]  ( .D(n280), .CK(clk), .Q(rs_id[1]), 
        .QN(n4402) );
  TBUF_X1 \ctrl_u/en_mul_id_tri  ( .A(\ctrl_u/n15 ), .EN(
        \ctrl_u/curr_mul_in_prog ), .Z(en_mul_id) );
  TBUF_X1 \ctrl_u/en_add_id_tri  ( .A(\ctrl_u/n11 ), .EN(
        \ctrl_u/curr_mul_in_prog ), .Z(en_add_id) );
  DFF_X1 \ctrl_u/curr_exe_reg[39]  ( .D(\ctrl_u/n422 ), .CK(clk), .Q(n4300), 
        .QN(\ctrl_u/curr_exe_39 ) );
  TBUF_X1 \ctrl_u/update_type_mem_tri[1]  ( .A(\ctrl_u/curr_mem_12 ), .EN(
        \ctrl_u/curr_ms ), .Z(dcache_update_type[1]) );
  TBUF_X1 \ctrl_u/update_type_mem_tri[0]  ( .A(\ctrl_u/curr_mem_11 ), .EN(
        \ctrl_u/curr_ms ), .Z(dcache_update_type[0]) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[25]  ( .D(n3048), .CK(clk), .Q(n4124), 
        .QN(n4211) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[63]  ( .D(n2819), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[63] ), .QN(n4583) );
  DFF_X1 \ctrl_u/curr_exe_reg[20]  ( .D(\ctrl_u/n441 ), .CK(clk), .Q(n4444), 
        .QN(\ctrl_u/curr_exe[20] ) );
  DFF_X1 \dp/ifs/pc/q_reg[25]  ( .D(n2532), .CK(clk), .Q(
        btb_cache_read_address[25]), .QN(n4599) );
  TBUF_X1 \ctrl_u/en_a_neg_id_tri  ( .A(1'b0), .EN(\ctrl_u/curr_mul_in_prog ), 
        .Z(en_a_neg_id) );
  TBUF_X1 \ctrl_u/en_a_neg_id_tri2  ( .A(n5158), .EN(n3933), .Z(en_a_neg_id)
         );
  DFF_X1 \ctrl_u/curr_exe_reg[28]  ( .D(\ctrl_u/n433 ), .CK(clk), .Q(n4236), 
        .QN(op_type_exe[0]) );
  DFF_X1 \ctrl_u/curr_id_reg[55]  ( .D(\ctrl_u/n509 ), .CK(clk), .Q(
        sign_ext_sel_id), .QN(n4448) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[61]  ( .D(n2821), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[61] ), .QN(n4452) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[63]  ( .D(n2883), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[63] ), .QN(n4493) );
  DFF_X1 \ctrl_u/curr_exe_reg[17]  ( .D(\ctrl_u/n444 ), .CK(clk), .Q(n4182), 
        .QN(\ctrl_u/curr_exe[17] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[10]  ( .D(\ctrl_u/n451 ), .CK(clk), .Q(n4450), 
        .QN(\ctrl_u/curr_exe[10] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[8]  ( .D(\ctrl_u/n453 ), .CK(clk), .Q(n4181), 
        .QN(\ctrl_u/curr_exe[8] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[7]  ( .D(\ctrl_u/n454 ), .CK(clk), .Q(n4180), 
        .QN(\ctrl_u/curr_exe[7] ) );
  TBUF_X1 \ctrl_u/shift_reg_id_tri  ( .A(1'b0), .EN(\ctrl_u/curr_mul_in_prog ), 
        .Z(shift_reg_id) );
  DFF_X1 \ctrl_u/curr_exe_reg[23]  ( .D(\ctrl_u/n438 ), .CK(clk), .Q(n4139), 
        .QN(alu_comp_sel[2]) );
  DFF_X1 \ctrl_u/curr_exe_reg[21]  ( .D(\ctrl_u/n440 ), .CK(clk), .Q(n4383), 
        .QN(alu_comp_sel[0]) );
  DFF_X1 \ctrl_u/curr_id_reg[53]  ( .D(\ctrl_u/n193 ), .CK(clk), .Q(n4357), 
        .QN(b_selector_id) );
  DFF_X1 \ctrl_u/curr_exe_reg[27]  ( .D(\ctrl_u/n434 ), .CK(clk), .Q(n4317), 
        .QN(op_sign_exe) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[17]  ( .D(n3056), .CK(clk), .Q(n4115), 
        .QN(n4205) );
  DFF_X1 \ctrl_u/curr_exe_reg[24]  ( .D(\ctrl_u/n437 ), .CK(clk), .Q(n4123), 
        .QN(cond_sel_exe[0]) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[38]  ( .D(n2844), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[38] ), .QN(n4474) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[37]  ( .D(n2845), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[37] ), .QN(n4473) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[24]  ( .D(n2922), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[24] ), .QN(n4284) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[58]  ( .D(n2824), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[58] ), .QN(n4442) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[24]  ( .D(n3049), .CK(clk), .Q(
        \dp/imm_id_exe_int[24] ), .QN(n4221) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[27]  ( .D(n2919), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[27] ), .QN(n4404) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[25]  ( .D(n2921), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[25] ), .QN(n4273) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[23]  ( .D(n2923), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[23] ), .QN(n4272) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[22]  ( .D(n2924), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[22] ), .QN(n4271) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[21]  ( .D(n2925), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[21] ), .QN(n4270) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[19]  ( .D(n2927), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[19] ), .QN(n4268) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[18]  ( .D(n2928), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[18] ), .QN(n4267) );
  TBUF_X1 \ctrl_u/en_imm_id_tri  ( .A(\ctrl_u/n27 ), .EN(
        \ctrl_u/curr_mul_in_prog ), .Z(en_imm_id) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[44]  ( .D(n2838), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[44] ), .QN(n4405) );
  DFF_X1 \ctrl_u/curr_exe_reg[15]  ( .D(\ctrl_u/n446 ), .CK(clk), .Q(n4167), 
        .QN(\ctrl_u/curr_exe[15] ) );
  DFF_X1 \ctrl_u/curr_exe_reg[25]  ( .D(\ctrl_u/n436 ), .CK(clk), .Q(n4126), 
        .QN(cond_sel_exe[1]) );
  DFF_X1 \ctrl_u/curr_exe_reg[26]  ( .D(\ctrl_u/n435 ), .CK(clk), .Q(n4494), 
        .QN(cond_sel_exe[2]) );
  DFF_X1 \ctrl_u/curr_exe_reg[35]  ( .D(\ctrl_u/n426 ), .CK(clk), .Q(n4445), 
        .QN(shift_type_exe[1]) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[20]  ( .D(n3053), .CK(clk), .QN(n4259)
         );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[18]  ( .D(n3055), .CK(clk), .QN(n4257)
         );
  TBUF_X1 \ctrl_u/en_b_id_tri  ( .A(\ctrl_u/n9 ), .EN(
        \ctrl_u/curr_mul_in_prog ), .Z(en_b_id) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[28]  ( .D(n2918), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[28] ), .QN(n4286) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[16]  ( .D(n3057), .CK(clk), .Q(
        \dp/imm_id_exe_int[16] ), .QN(n4219) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[56]  ( .D(n2826), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[56] ), .QN(n4387) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[51]  ( .D(n2831), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[51] ), .QN(n6620) );
  TBUF_X1 \ctrl_u/en_shift_id_tri  ( .A(\ctrl_u/n13 ), .EN(
        \ctrl_u/curr_mul_in_prog ), .Z(en_shift_id) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[33]  ( .D(n2849), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[33] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[48]  ( .D(n2898), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[48] ) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[21]  ( .D(n279), .CK(clk), .Q(rs_id[0]), 
        .QN(n4083) );
  DFF_X1 \dp/ex_mem_regs/alu_out_low_reg/q_reg[4]  ( .D(n2649), .CK(clk), .Q(
        \dp/mul_feedback_exe_mem_int[4] ), .QN(n4071) );
  TBUF_X1 \ctrl_u/en_npc_id_tri  ( .A(\ctrl_u/n25 ), .EN(
        \ctrl_u/curr_mul_in_prog ), .Z(en_npc_id) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[52]  ( .D(n2830), .CK(clk), .Q(
        \dp/a_neg_mult_id_exe_int[52] ), .QN(n4380) );
  DFF_X1 \ctrl_u/curr_exe_reg[34]  ( .D(\ctrl_u/n427 ), .CK(clk), .Q(n4378), 
        .QN(shift_type_exe[0]) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[23]  ( .D(n281), .CK(clk), .Q(rs_id[2]), 
        .QN(n4370) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[19]  ( .D(n277), .CK(clk), .Q(rt_id[3]), 
        .QN(n4212) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[18]  ( .D(n276), .CK(clk), .Q(rt_id[2]), 
        .QN(n4365) );
  TBUF_X1 \ctrl_u/en_rd_id_tri  ( .A(\ctrl_u/n23 ), .EN(
        \ctrl_u/curr_mul_in_prog ), .Z(en_rd_id) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[25]  ( .D(n283), .CK(clk), .Q(rs_id[4]), 
        .QN(n4360) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[20]  ( .D(n278), .CK(clk), .Q(rt_id[4]), 
        .QN(n4359) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[16]  ( .D(n274), .CK(clk), .Q(rt_id[0]), 
        .QN(n7172) );
  DFF_X1 \dp/if_id_regs/ir_reg/q_reg[24]  ( .D(n282), .CK(clk), .Q(rs_id[3]), 
        .QN(n4366) );
  TBUF_X1 \ctrl_u/en_shift_reg_id_tri  ( .A(\ctrl_u/n21 ), .EN(
        \ctrl_u/curr_mul_in_prog ), .Z(en_shift_reg_id) );
  NAND2_X1 \intadd_1/U29  ( .A1(\intadd_1/A[23] ), .A2(\intadd_1/B[23] ), .ZN(
        \intadd_1/n45 ) );
  NAND2_X1 \intadd_1/U19  ( .A1(\intadd_1/A[24] ), .A2(\intadd_1/B[24] ), .ZN(
        \intadd_1/n38 ) );
  NAND2_X1 \intadd_1/U132  ( .A1(\intadd_1/n188 ), .A2(\intadd_1/n115 ), .ZN(
        \intadd_1/n15 ) );
  XOR2_X1 \intadd_1/U213  ( .A(\intadd_1/n169 ), .B(\intadd_1/n25 ), .Z(
        \intadd_1/SUM[1] ) );
  NAND2_X1 \intadd_1/U222  ( .A1(\intadd_1/n199 ), .A2(\intadd_1/n172 ), .ZN(
        \intadd_1/n26 ) );
  NAND2_X1 \intadd_1/U200  ( .A1(\intadd_1/n196 ), .A2(\intadd_1/n159 ), .ZN(
        \intadd_1/n23 ) );
  XNOR2_X1 \intadd_1/U196  ( .A(\intadd_1/n160 ), .B(\intadd_1/n23 ), .ZN(
        \intadd_1/SUM[3] ) );
  NAND2_X1 \intadd_1/U209  ( .A1(n4045), .A2(\intadd_1/n165 ), .ZN(
        \intadd_1/n24 ) );
  XNOR2_X1 \intadd_1/U204  ( .A(\intadd_1/n166 ), .B(\intadd_1/n24 ), .ZN(
        \intadd_1/SUM[2] ) );
  NAND2_X1 \intadd_1/U178  ( .A1(\intadd_1/n193 ), .A2(\intadd_1/n146 ), .ZN(
        \intadd_1/n20 ) );
  NAND2_X1 \intadd_1/U114  ( .A1(\intadd_1/n186 ), .A2(\intadd_1/n103 ), .ZN(
        \intadd_1/n13 ) );
  NAND2_X1 \intadd_1/U71  ( .A1(\intadd_1/n181 ), .A2(\intadd_1/n75 ), .ZN(
        \intadd_1/n8 ) );
  AOI21_X1 \intadd_1/U111  ( .B1(\intadd_1/n104 ), .B2(\intadd_1/n186 ), .A(
        \intadd_1/n101 ), .ZN(\intadd_1/n99 ) );
  NAND2_X1 \intadd_1/U106  ( .A1(\intadd_1/n185 ), .A2(\intadd_1/n98 ), .ZN(
        \intadd_1/n12 ) );
  XOR2_X1 \intadd_1/U97  ( .A(\intadd_1/n99 ), .B(\intadd_1/n12 ), .Z(
        \intadd_1/SUM[14] ) );
  NAND2_X1 \intadd_1/U161  ( .A1(\intadd_1/n191 ), .A2(\intadd_1/n135 ), .ZN(
        \intadd_1/n18 ) );
  XNOR2_X1 \intadd_1/U155  ( .A(\intadd_1/n136 ), .B(\intadd_1/n18 ), .ZN(
        \intadd_1/SUM[8] ) );
  NAND2_X1 \intadd_1/U38  ( .A1(\intadd_1/n177 ), .A2(\intadd_1/n54 ), .ZN(
        \intadd_1/n4 ) );
  AOI21_X1 \intadd_1/U129  ( .B1(\intadd_1/n117 ), .B2(\intadd_1/n188 ), .A(
        \intadd_1/n113 ), .ZN(\intadd_1/n111 ) );
  NAND2_X1 \intadd_1/U124  ( .A1(n3914), .A2(\intadd_1/n110 ), .ZN(
        \intadd_1/n14 ) );
  XOR2_X1 \intadd_1/U118  ( .A(\intadd_1/n111 ), .B(\intadd_1/n14 ), .Z(
        \intadd_1/SUM[12] ) );
  NAND2_X1 \intadd_1/U52  ( .A1(\intadd_1/n179 ), .A2(\intadd_1/n62 ), .ZN(
        \intadd_1/n6 ) );
  XNOR2_X1 \intadd_1/U48  ( .A(\intadd_1/n63 ), .B(\intadd_1/n6 ), .ZN(
        \intadd_1/SUM[20] ) );
  HA_X1 \add_x_20/U27  ( .A(\add_x_20/n27 ), .B(btb_cache_read_address[3]), 
        .CO(\add_x_20/n26 ), .S(\dp/pc_plus4_out_if_int[3] ) );
  HA_X1 \add_x_20/U26  ( .A(\add_x_20/n26 ), .B(btb_cache_read_address[4]), 
        .CO(\add_x_20/n25 ), .S(\dp/pc_plus4_out_if_int[4] ) );
  HA_X1 \add_x_20/U25  ( .A(\add_x_20/n25 ), .B(btb_cache_read_address[5]), 
        .CO(\add_x_20/n24 ), .S(\dp/pc_plus4_out_if_int[5] ) );
  HA_X1 \add_x_20/U24  ( .A(\add_x_20/n24 ), .B(btb_cache_read_address[6]), 
        .CO(\add_x_20/n23 ), .S(\dp/pc_plus4_out_if_int[6] ) );
  HA_X1 \add_x_20/U23  ( .A(\add_x_20/n23 ), .B(btb_cache_read_address[7]), 
        .CO(\add_x_20/n22 ), .S(\dp/pc_plus4_out_if_int[7] ) );
  HA_X1 \add_x_20/U22  ( .A(\add_x_20/n22 ), .B(btb_cache_read_address[8]), 
        .CO(\add_x_20/n21 ), .S(\dp/pc_plus4_out_if_int[8] ) );
  HA_X1 \add_x_20/U21  ( .A(\add_x_20/n21 ), .B(btb_cache_read_address[9]), 
        .CO(\add_x_20/n20 ), .S(\dp/pc_plus4_out_if_int[9] ) );
  HA_X1 \add_x_20/U20  ( .A(\add_x_20/n20 ), .B(btb_cache_read_address[10]), 
        .CO(\add_x_20/n19 ), .S(\dp/pc_plus4_out_if_int[10] ) );
  HA_X1 \add_x_20/U19  ( .A(\add_x_20/n19 ), .B(btb_cache_read_address[11]), 
        .CO(\add_x_20/n18 ), .S(\dp/pc_plus4_out_if_int[11] ) );
  HA_X1 \add_x_20/U18  ( .A(\add_x_20/n18 ), .B(btb_cache_read_address[12]), 
        .CO(\add_x_20/n17 ), .S(\dp/pc_plus4_out_if_int[12] ) );
  HA_X1 \add_x_20/U17  ( .A(\add_x_20/n17 ), .B(btb_cache_read_address[13]), 
        .CO(\add_x_20/n16 ), .S(\dp/pc_plus4_out_if_int[13] ) );
  HA_X1 \add_x_20/U16  ( .A(\add_x_20/n16 ), .B(btb_cache_read_address[14]), 
        .CO(\add_x_20/n15 ), .S(\dp/pc_plus4_out_if_int[14] ) );
  HA_X1 \add_x_20/U15  ( .A(\add_x_20/n15 ), .B(btb_cache_read_address[15]), 
        .CO(\add_x_20/n14 ), .S(\dp/pc_plus4_out_if_int[15] ) );
  HA_X1 \add_x_20/U14  ( .A(\add_x_20/n14 ), .B(btb_cache_read_address[16]), 
        .CO(\add_x_20/n13 ), .S(\dp/pc_plus4_out_if_int[16] ) );
  HA_X1 \add_x_20/U13  ( .A(\add_x_20/n13 ), .B(btb_cache_read_address[17]), 
        .CO(\add_x_20/n12 ), .S(\dp/pc_plus4_out_if_int[17] ) );
  HA_X1 \add_x_20/U12  ( .A(\add_x_20/n12 ), .B(btb_cache_read_address[18]), 
        .CO(\add_x_20/n11 ), .S(\dp/pc_plus4_out_if_int[18] ) );
  HA_X1 \add_x_20/U11  ( .A(\add_x_20/n11 ), .B(btb_cache_read_address[19]), 
        .CO(\add_x_20/n10 ), .S(\dp/pc_plus4_out_if_int[19] ) );
  HA_X1 \add_x_20/U10  ( .A(\add_x_20/n10 ), .B(btb_cache_read_address[20]), 
        .CO(\add_x_20/n9 ), .S(\dp/pc_plus4_out_if_int[20] ) );
  HA_X1 \add_x_20/U9  ( .A(\add_x_20/n9 ), .B(btb_cache_read_address[21]), 
        .CO(\add_x_20/n8 ), .S(\dp/pc_plus4_out_if_int[21] ) );
  HA_X1 \add_x_20/U8  ( .A(\add_x_20/n8 ), .B(btb_cache_read_address[22]), 
        .CO(\add_x_20/n7 ), .S(\dp/pc_plus4_out_if_int[22] ) );
  HA_X1 \add_x_20/U7  ( .A(\add_x_20/n7 ), .B(btb_cache_read_address[23]), 
        .CO(\add_x_20/n6 ), .S(\dp/pc_plus4_out_if_int[23] ) );
  HA_X1 \add_x_20/U6  ( .A(\add_x_20/n6 ), .B(btb_cache_read_address[24]), 
        .CO(\add_x_20/n5 ), .S(\dp/pc_plus4_out_if_int[24] ) );
  HA_X1 \add_x_20/U5  ( .A(\add_x_20/n5 ), .B(btb_cache_read_address[25]), 
        .CO(\add_x_20/n4 ), .S(\dp/pc_plus4_out_if_int[25] ) );
  HA_X1 \add_x_20/U4  ( .A(\add_x_20/n4 ), .B(btb_cache_read_address[26]), 
        .CO(\add_x_20/n3 ), .S(\dp/pc_plus4_out_if_int[26] ) );
  HA_X1 \add_x_20/U3  ( .A(\add_x_20/n3 ), .B(btb_cache_read_address[27]), 
        .CO(\add_x_20/n2 ), .S(\dp/pc_plus4_out_if_int[27] ) );
  DFF_X1 \dp/mem_wb_regs/rd_reg/q_reg[1]  ( .D(n1598), .CK(clk), .Q(n4005), 
        .QN(n7537) );
  DFF_X2 \ctrl_u/curr_id_reg[54]  ( .D(\ctrl_u/n510 ), .CK(clk), .Q(n4136), 
        .QN(n4358) );
  DFF_X1 \dp/mem_wb_regs/rd_reg/q_reg[4]  ( .D(n1688), .CK(clk), .QN(n7534) );
  DFF_X1 \dp/mem_wb_regs/rd_reg/q_reg[3]  ( .D(n1594), .CK(clk), .QN(n7535) );
  DFF_X1 \dp/mem_wb_regs/rd_reg/q_reg[2]  ( .D(n1597), .CK(clk), .QN(n7536) );
  DFF_X1 \dp/mem_wb_regs/rd_reg/q_reg[0]  ( .D(n1599), .CK(clk), .QN(n7538) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[7]  ( .D(n1680), .CK(clk), .QN(
        \dp/cache_data_mem_wb_int[7] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[6]  ( .D(n1681), .CK(clk), .QN(
        \dp/cache_data_mem_wb_int[6] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[5]  ( .D(n1682), .CK(clk), .QN(
        \dp/cache_data_mem_wb_int[5] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[4]  ( .D(n1683), .CK(clk), .QN(
        \dp/cache_data_mem_wb_int[4] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[3]  ( .D(n1684), .CK(clk), .QN(
        \dp/cache_data_mem_wb_int[3] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[2]  ( .D(n1685), .CK(clk), .QN(
        \dp/cache_data_mem_wb_int[2] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[1]  ( .D(n1686), .CK(clk), .QN(
        \dp/cache_data_mem_wb_int[1] ) );
  DFF_X1 \dp/mem_wb_regs/cache_data_reg/q_reg[0]  ( .D(n1687), .CK(clk), .QN(
        \dp/cache_data_mem_wb_int[0] ) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[17]  ( .D(n1459), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[17] ) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[19]  ( .D(n1457), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[19] ) );
  DFF_X1 \dp/id_exe_regs/npc_reg/q_reg[9]  ( .D(n3001), .CK(clk), .QN(n4217)
         );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[27]  ( .D(n3046), .CK(clk), .QN(n4398)
         );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[20]  ( .D(n1456), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[20] ) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[18]  ( .D(n1458), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[18] ) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[16]  ( .D(n1460), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[16] ) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[21]  ( .D(n1455), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[21] ) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[15]  ( .D(n1461), .CK(clk), .QN(
        \dp/a_neg_mult_id_exe_int[15] ) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[1]  ( .D(n1143), .CK(clk), .QN(
        \dp/op_b_id_ex_int[1] ) );
  DFF_X1 \dp/id_exe_regs/b_reg/q_reg[0]  ( .D(n1144), .CK(clk), .QN(
        \dp/op_b_id_ex_int[0] ) );
  DFF_X1 \dp/id_exe_regs/b_shift_reg/q_reg[4]  ( .D(n2717), .CK(clk), .QN(
        n4260) );
  DFF_X1 \dp/id_exe_regs/b_shift_reg/q_reg[1]  ( .D(n2720), .CK(clk), .QN(
        n4263) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[29]  ( .D(n2949), .CK(clk), .QN(
        n642) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[25]  ( .D(n2953), .CK(clk), .QN(
        n638) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[21]  ( .D(n2957), .CK(clk), .QN(
        n634) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[17]  ( .D(n2961), .CK(clk), .QN(
        n630) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[14]  ( .D(n2964), .CK(clk), .QN(
        n627) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[13]  ( .D(n2965), .CK(clk), .QN(
        n626) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[5]  ( .D(n2973), .CK(clk), .QN(n618) );
  DFF_X1 \dp/id_exe_regs/b_shift_reg/q_reg[3]  ( .D(n2718), .CK(clk), .QN(
        n4261) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[31]  ( .D(n2947), .CK(clk), .QN(
        n644) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[26]  ( .D(n2952), .CK(clk), .QN(
        n639) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[22]  ( .D(n2956), .CK(clk), .QN(
        n635) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[10]  ( .D(n2968), .CK(clk), .QN(
        n623) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[27]  ( .D(n2951), .CK(clk), .QN(
        n640) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[24]  ( .D(n2954), .CK(clk), .QN(
        n637) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[23]  ( .D(n2955), .CK(clk), .QN(
        n636) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[20]  ( .D(n2958), .CK(clk), .QN(
        n633) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[19]  ( .D(n2959), .CK(clk), .QN(
        n632) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[16]  ( .D(n2962), .CK(clk), .QN(
        n629) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[15]  ( .D(n2963), .CK(clk), .QN(
        n628) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[12]  ( .D(n2966), .CK(clk), .QN(
        n625) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[11]  ( .D(n2967), .CK(clk), .QN(
        n624) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[8]  ( .D(n2970), .CK(clk), .QN(n621) );
  DFF_X1 \dp/id_exe_regs/b_shift_reg/q_reg[2]  ( .D(n2719), .CK(clk), .QN(
        n4262) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[30]  ( .D(n2948), .CK(clk), .QN(
        n643) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[18]  ( .D(n2960), .CK(clk), .QN(
        n631) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[9]  ( .D(n2969), .CK(clk), .QN(n622) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[6]  ( .D(n2972), .CK(clk), .QN(n619) );
  DFF_X1 \dp/id_exe_regs/b_shift_reg/q_reg[0]  ( .D(n2721), .CK(clk), .QN(
        n4264) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[2]  ( .D(n2976), .CK(clk), .QN(n615) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[9]  ( .D(n259), .CK(clk), .QN(
        \intadd_2/A[6] ) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[19]  ( .D(n3054), .CK(clk), .QN(n4258)
         );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[28]  ( .D(n2950), .CK(clk), .QN(
        n641) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[7]  ( .D(n2971), .CK(clk), .QN(n620) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[4]  ( .D(n2974), .CK(clk), .QN(n617) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[3]  ( .D(n2975), .CK(clk), .QN(n616) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[1]  ( .D(n2977), .CK(clk), .QN(n614) );
  DFF_X1 \dp/id_exe_regs/a_shift_reg/q_reg[0]  ( .D(n2978), .CK(clk), .QN(n613) );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[28]  ( .D(n3045), .CK(clk), .QN(n4399)
         );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[29]  ( .D(n3044), .CK(clk), .QN(n4400)
         );
  DFF_X1 \dp/id_exe_regs/imm_reg/q_reg[26]  ( .D(n3047), .CK(clk), .QN(n4397)
         );
  DFF_X1 \ctrl_u/curr_mul_end_mem_reg  ( .D(\ctrl_u/n560 ), .CK(clk), .Q(
        \ctrl_u/curr_mul_end_mem ) );
  DFF_X1 \ctrl_u/curr_id_reg[22]  ( .D(\ctrl_u/n536 ), .CK(clk), .Q(
        \ctrl_u/curr_id[22] ) );
  DFF_X1 \ctrl_u/curr_id_reg[0]  ( .D(\ctrl_u/n553 ), .CK(clk), .Q(
        \ctrl_u/curr_id[0] ), .QN(n5566) );
  DFF_X1 \ctrl_u/curr_id_reg[39]  ( .D(\ctrl_u/n523 ), .CK(clk), .Q(
        \ctrl_u/curr_id[39] ) );
  DFF_X1 \ctrl_u/curr_id_reg[12]  ( .D(\ctrl_u/n544 ), .CK(clk), .Q(
        \ctrl_u/curr_id[12] ), .QN(n5555) );
  DFF_X1 \ctrl_u/curr_id_reg[60]  ( .D(\ctrl_u/n506 ), .CK(clk), .Q(
        rp1_out_sel_id[1]), .QN(n5485) );
  DFF_X1 \ctrl_u/curr_id_reg[59]  ( .D(\ctrl_u/n507 ), .CK(clk), .Q(
        rp1_out_sel_id[0]), .QN(n5487) );
  DFF_X1 \ctrl_u/curr_id_reg[28]  ( .D(\ctrl_u/n531 ), .CK(clk), .Q(
        \ctrl_u/curr_id[28] ) );
  DFF_X2 \ctrl_u/curr_wb_reg[1]  ( .D(\ctrl_u/n484 ), .CK(clk), .Q(n4336), 
        .QN(n5228) );
  DFF_X1 \dp/ifs/pc/q_reg[28]  ( .D(n2529), .CK(clk), .Q(
        btb_cache_read_address[28]), .QN(n3869) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[0]  ( .D(n2946), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[0] ), .QN(n4369) );
  DFF_X1 \ctrl_u/curr_mem_reg[3]  ( .D(\ctrl_u/n477 ), .CK(clk), .Q(n4265), 
        .QN(\ctrl_u/curr_mem[3] ) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[1]  ( .D(n2945), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[1] ), .QN(n4230) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[5]  ( .D(n2941), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[5] ), .QN(n4223) );
  DFF_X1 \dp/id_exe_regs/a_mult_reg/q_reg[4]  ( .D(n2942), .CK(clk), .Q(
        \dp/a_mult_id_exe_int[4] ), .QN(n4108) );
  DFF_X1 \dp/id_exe_regs/a_neg_mult_reg/q_reg[5]  ( .D(n1471), .CK(clk), .Q(
        n4104), .QN(\dp/a_neg_mult_id_exe_int[5] ) );
  DFF_X1 \dp/ex_mem_regs/alu_out_high_reg/q_reg[22]  ( .D(n2796), .CK(clk), 
        .Q(\dp/mul_feedback_exe_mem_int[54] ), .QN(n4195) );
  OAI33_X1 U3011 ( .A1(1'b0), .A2(n3641), .A3(1'b0), .B1(n5099), .B2(n4785), 
        .B3(n4787), .ZN(n4781) );
  NOR2_X1 U3012 ( .A1(\intadd_1/A[14] ), .A2(\intadd_1/B[14] ), .ZN(
        \intadd_1/n97 ) );
  INV_X1 U3013 ( .A(n5330), .ZN(n3950) );
  BUF_X1 U3014 ( .A(n5168), .Z(n3899) );
  BUF_X2 U3015 ( .A(n5141), .Z(n5136) );
  AND4_X1 U3016 ( .A1(n5706), .A2(n5707), .A3(n5705), .A4(n5704), .ZN(n3911)
         );
  INV_X1 U3017 ( .A(n3911), .ZN(n5855) );
  INV_X1 U3018 ( .A(n6322), .ZN(n3951) );
  BUF_X2 U3019 ( .A(n7253), .Z(n5175) );
  AND2_X1 U3020 ( .A1(n5816), .A2(n5814), .ZN(n5842) );
  OR2_X1 U3021 ( .A1(n5680), .A2(n5679), .ZN(n5150) );
  NAND2_X1 U3022 ( .A1(n5751), .A2(log_type_exe[2]), .ZN(n7080) );
  INV_X1 U3023 ( .A(n5027), .ZN(n3948) );
  INV_X1 U3024 ( .A(n5581), .ZN(n3941) );
  CLKBUF_X3 U3025 ( .A(n7104), .Z(n3879) );
  AOI21_X1 U3026 ( .B1(n6111), .B2(n7076), .A(n6110), .ZN(n6416) );
  BUF_X2 U3027 ( .A(n6756), .Z(n4055) );
  BUF_X2 U3028 ( .A(n4224), .Z(n3897) );
  BUF_X2 U3029 ( .A(n4224), .Z(n3896) );
  BUF_X2 U3030 ( .A(n4224), .Z(n3898) );
  BUF_X2 U3031 ( .A(n7036), .Z(n3881) );
  BUF_X2 U3032 ( .A(n7036), .Z(n3880) );
  NAND2_X1 U3033 ( .A1(n3989), .A2(n3952), .ZN(n5812) );
  AOI22_X1 U3034 ( .A1(n5154), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[51] ), 
        .B1(n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[52] ), .ZN(n3268) );
  NAND2_X1 U3035 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[52] ), .A2(n5188), 
        .ZN(n3269) );
  OAI21_X1 U3036 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[52] ), .A(n3269), 
        .ZN(n3270) );
  AOI21_X1 U3037 ( .B1(n5189), .B2(\dp/exs/alu_unit/mult/a_shiftn[51] ), .A(
        n3270), .ZN(n3271) );
  NAND2_X1 U3038 ( .A1(n3268), .A2(n3271), .ZN(n6277) );
  NOR2_X1 U3039 ( .A1(n5230), .A2(n380), .ZN(n3272) );
  AOI21_X1 U3040 ( .B1(\dp/ids/rp1[22] ), .B2(n4136), .A(n3272), .ZN(n6811) );
  INV_X1 U3041 ( .A(n7056), .ZN(n3273) );
  NAND2_X1 U3042 ( .A1(\dp/a_mult_id_exe_int[17] ), .A2(n3878), .ZN(n3274) );
  OAI21_X1 U3043 ( .B1(n3273), .B2(n6835), .A(n3274), .ZN(n2929) );
  AOI22_X1 U3044 ( .A1(n5184), .A2(\dp/a_neg_mult_id_exe_int[33] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[33] ), .ZN(n3275) );
  AOI22_X1 U3045 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[32] ), .B1(
        \dp/mul_feedback_exe_mem_int[33] ), .B2(n5186), .ZN(n3276) );
  NAND2_X1 U3046 ( .A1(n3275), .A2(n3276), .ZN(n6197) );
  AOI22_X1 U3047 ( .A1(n3945), .A2(\dp/exs/alu_unit/mult/a_shiftn[56] ), .B1(
        n5189), .B2(\dp/exs/alu_unit/mult/a_shiftn[55] ), .ZN(n3277) );
  NAND2_X1 U3048 ( .A1(n3946), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[56] ), 
        .ZN(n3278) );
  OAI21_X1 U3049 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[56] ), .A(n3278), 
        .ZN(n3279) );
  AOI21_X1 U3050 ( .B1(n5154), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[55] ), 
        .A(n3279), .ZN(n3280) );
  NAND2_X1 U3051 ( .A1(n3277), .A2(n3280), .ZN(n6289) );
  AOI22_X1 U3052 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/a_shiftn[16] ), .B1(
        n3946), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[17] ), .ZN(n3281) );
  NAND2_X1 U3053 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[17] ), .A2(n3945), .ZN(
        n3282) );
  OAI21_X1 U3054 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[17] ), .A(n3282), 
        .ZN(n3283) );
  AOI21_X1 U3055 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[16] ), 
        .A(n3283), .ZN(n3284) );
  NAND2_X1 U3056 ( .A1(n3281), .A2(n3284), .ZN(n5956) );
  NOR2_X1 U3057 ( .A1(n5230), .A2(n379), .ZN(n3285) );
  AOI21_X1 U3058 ( .B1(\dp/ids/rp1[21] ), .B2(n4136), .A(n3285), .ZN(n6816) );
  AOI22_X1 U3059 ( .A1(\dp/a_neg_mult_id_exe_int[19] ), .A2(n7098), .B1(n6429), 
        .B2(n7097), .ZN(n1457) );
  INV_X1 U3060 ( .A(n5200), .ZN(n3286) );
  NAND2_X1 U3061 ( .A1(\dp/a_mult_id_exe_int[16] ), .A2(n3876), .ZN(n3287) );
  OAI21_X1 U3062 ( .B1(n3286), .B2(n6838), .A(n3287), .ZN(n2930) );
  AOI22_X1 U3063 ( .A1(n3943), .A2(\dp/a_neg_mult_id_exe_int[34] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[35] ), .ZN(n3288) );
  AOI22_X1 U3064 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[35] ), .B1(
        \dp/mul_feedback_exe_mem_int[35] ), .B2(n5186), .ZN(n3289) );
  NAND2_X1 U3065 ( .A1(n3288), .A2(n3289), .ZN(n6201) );
  AOI22_X1 U3066 ( .A1(n5184), .A2(\dp/a_neg_mult_id_exe_int[39] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[39] ), .ZN(n3290) );
  AOI22_X1 U3067 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[38] ), .B1(
        \dp/mul_feedback_exe_mem_int[39] ), .B2(n5186), .ZN(n3291) );
  NAND2_X1 U3068 ( .A1(n3290), .A2(n3291), .ZN(n6218) );
  AOI22_X1 U3069 ( .A1(n5188), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[54] ), 
        .B1(n5189), .B2(\dp/exs/alu_unit/mult/a_shiftn[53] ), .ZN(n3292) );
  NAND2_X1 U3070 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[53] ), .A2(n6326), 
        .ZN(n3293) );
  OAI21_X1 U3071 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[54] ), .A(n3293), 
        .ZN(n3294) );
  AOI21_X1 U3072 ( .B1(n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[54] ), .A(
        n3294), .ZN(n3295) );
  NAND2_X1 U3073 ( .A1(n3292), .A2(n3295), .ZN(n6284) );
  AOI22_X1 U3074 ( .A1(n5154), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[56] ), 
        .B1(n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[57] ), .ZN(n3296) );
  NAND2_X1 U3075 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[57] ), .A2(n3946), 
        .ZN(n3297) );
  OAI21_X1 U3076 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[57] ), .A(n3297), 
        .ZN(n3298) );
  AOI21_X1 U3077 ( .B1(n5189), .B2(\dp/exs/alu_unit/mult/a_shiftn[56] ), .A(
        n3298), .ZN(n3299) );
  NAND2_X1 U3078 ( .A1(n3296), .A2(n3299), .ZN(n6291) );
  NOR2_X1 U3079 ( .A1(n7080), .A2(n6163), .ZN(n3300) );
  AOI21_X1 U3080 ( .B1(n6159), .B2(n6160), .A(n3300), .ZN(n3301) );
  XNOR2_X1 U3081 ( .A(n6309), .B(n6156), .ZN(n3302) );
  AOI22_X1 U3082 ( .A1(n3954), .A2(\dp/exs/alu_unit/shifter_out[31] ), .B1(
        n7076), .B2(n3302), .ZN(n3303) );
  OAI211_X1 U3083 ( .C1(n6164), .C2(n7066), .A(n3301), .B(n3303), .ZN(n6410)
         );
  NOR2_X1 U3084 ( .A1(n5230), .A2(n378), .ZN(n3304) );
  AOI21_X1 U3085 ( .B1(\dp/ids/rp1[20] ), .B2(n4136), .A(n3304), .ZN(n6821) );
  AOI22_X1 U3086 ( .A1(\dp/a_neg_mult_id_exe_int[17] ), .A2(n7098), .B1(n4910), 
        .B2(n7097), .ZN(n1459) );
  INV_X1 U3087 ( .A(n5201), .ZN(n3305) );
  NAND2_X1 U3088 ( .A1(\dp/a_mult_id_exe_int[15] ), .A2(n3877), .ZN(n3306) );
  OAI21_X1 U3089 ( .B1(n3305), .B2(n6841), .A(n3306), .ZN(n2931) );
  AOI22_X1 U3090 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/a_shiftn[29] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[30] ), .ZN(n3307) );
  NAND2_X1 U3091 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[29] ), .A2(n6326), 
        .ZN(n3308) );
  OAI21_X1 U3092 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[30] ), .A(n3308), 
        .ZN(n3309) );
  AOI21_X1 U3093 ( .B1(n3946), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[30] ), 
        .A(n3309), .ZN(n3310) );
  NAND2_X1 U3094 ( .A1(n3307), .A2(n3310), .ZN(n6139) );
  AOI22_X1 U3095 ( .A1(n5184), .A2(\dp/a_neg_mult_id_exe_int[43] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[43] ), .ZN(n3311) );
  AOI22_X1 U3096 ( .A1(n3943), .A2(\dp/a_neg_mult_id_exe_int[42] ), .B1(
        \dp/mul_feedback_exe_mem_int[43] ), .B2(n5186), .ZN(n3312) );
  NAND2_X1 U3097 ( .A1(n3311), .A2(n3312), .ZN(n6244) );
  AOI22_X1 U3098 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/a_shiftn[59] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[60] ), .ZN(n3313) );
  NAND2_X1 U3099 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[59] ), .A2(n5154), 
        .ZN(n3314) );
  OAI21_X1 U3100 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[60] ), .A(n3314), 
        .ZN(n3315) );
  AOI21_X1 U3101 ( .B1(n3946), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[60] ), 
        .A(n3315), .ZN(n3316) );
  NAND2_X1 U3102 ( .A1(n3313), .A2(n3316), .ZN(n6300) );
  AOI22_X1 U3103 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/a_shiftn[14] ), .B1(
        n3946), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[15] ), .ZN(n3317) );
  NAND2_X1 U3104 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[15] ), .A2(n3945), .ZN(
        n3318) );
  OAI21_X1 U3105 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[15] ), .A(n3318), 
        .ZN(n3319) );
  AOI21_X1 U3106 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[14] ), 
        .A(n3319), .ZN(n3320) );
  NAND2_X1 U3107 ( .A1(n3317), .A2(n3320), .ZN(n5943) );
  AOI22_X1 U3108 ( .A1(n6326), .A2(\dp/exs/alu_unit/mult/neg_ax2_shiftn[12] ), 
        .B1(n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[12] ), .ZN(n3321) );
  NAND2_X1 U3109 ( .A1(\dp/exs/alu_unit/mult/ax2_shiftn[12] ), .A2(n5189), 
        .ZN(n3322) );
  OAI21_X1 U3110 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[12] ), .A(n3322), 
        .ZN(n3323) );
  AOI21_X1 U3111 ( .B1(n3946), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[12] ), 
        .A(n3323), .ZN(n3324) );
  NAND2_X1 U3112 ( .A1(n3321), .A2(n3324), .ZN(n5925) );
  AOI22_X1 U3113 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/ax2_shiftn[9] ), .B1(
        n5188), .B2(\dp/exs/alu_unit/mult/neg_ax2_shiftn[10] ), .ZN(n3325) );
  NAND2_X1 U3114 ( .A1(\dp/exs/alu_unit/mult/ax2_shiftn[10] ), .A2(n3945), 
        .ZN(n3326) );
  OAI21_X1 U3115 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[9] ), .A(n3326), .ZN(
        n3327) );
  AOI21_X1 U3116 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_ax2_shiftn[9] ), 
        .A(n3327), .ZN(n3328) );
  NAND2_X1 U3117 ( .A1(n3325), .A2(n3328), .ZN(n5909) );
  XNOR2_X1 U3118 ( .A(n6119), .B(n6141), .ZN(n3329) );
  XNOR2_X1 U3119 ( .A(n3329), .B(n6118), .ZN(n3330) );
  INV_X1 U3120 ( .A(n6113), .ZN(n3331) );
  AOI221_X1 U3121 ( .B1(n7069), .B2(n3331), .C1(n7080), .C2(n6113), .A(
        \intadd_1/B[28] ), .ZN(n3332) );
  AOI21_X1 U3122 ( .B1(n3954), .B2(\dp/exs/alu_unit/shifter_out[29] ), .A(
        n3332), .ZN(n3333) );
  NAND3_X1 U3123 ( .A1(\intadd_1/B[28] ), .A2(n3952), .A3(n3331), .ZN(n3334)
         );
  OAI211_X1 U3124 ( .C1(n3864), .C2(n7066), .A(n3333), .B(n3334), .ZN(n3335)
         );
  AOI21_X1 U3125 ( .B1(n3330), .B2(n7076), .A(n3335), .ZN(n6414) );
  NOR2_X1 U3126 ( .A1(n5230), .A2(n369), .ZN(n3336) );
  AOI21_X1 U3127 ( .B1(\dp/ids/rp1[11] ), .B2(n4136), .A(n3336), .ZN(n6851) );
  NAND2_X1 U3128 ( .A1(n5644), .A2(instr_if[28]), .ZN(n3337) );
  AOI22_X1 U3129 ( .A1(n5645), .A2(n5646), .B1(n5647), .B2(n3337), .ZN(n3338)
         );
  AOI221_X1 U3130 ( .B1(n5650), .B2(n5648), .C1(n5649), .C2(n5648), .A(n5643), 
        .ZN(n3339) );
  NAND3_X1 U3131 ( .A1(n5651), .A2(n3338), .A3(n3339), .ZN(n3340) );
  OAI22_X1 U3132 ( .A1(b_selector_id), .A2(n5652), .B1(n3927), .B2(n3340), 
        .ZN(\ctrl_u/n193 ) );
  AOI22_X1 U3133 ( .A1(\dp/a_neg_mult_id_exe_int[25] ), .A2(n5126), .B1(n4895), 
        .B2(n7097), .ZN(n1451) );
  INV_X1 U3134 ( .A(n5202), .ZN(n3341) );
  NAND2_X1 U3135 ( .A1(\dp/a_mult_id_exe_int[14] ), .A2(n3877), .ZN(n3342) );
  OAI21_X1 U3136 ( .B1(n3341), .B2(n6844), .A(n3342), .ZN(n2932) );
  AND3_X1 U3137 ( .A1(n4726), .A2(n5096), .A3(n3961), .ZN(n5330) );
  AOI22_X1 U3138 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/a_shiftn[34] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[35] ), .ZN(n3343) );
  NAND2_X1 U3139 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[34] ), .A2(n6326), 
        .ZN(n3344) );
  OAI21_X1 U3140 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[35] ), .A(n3344), 
        .ZN(n3345) );
  AOI21_X1 U3141 ( .B1(n3946), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[35] ), 
        .A(n3345), .ZN(n3346) );
  NAND2_X1 U3142 ( .A1(n3343), .A2(n3346), .ZN(n6202) );
  AOI22_X1 U3143 ( .A1(n5184), .A2(\dp/a_neg_mult_id_exe_int[40] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[40] ), .ZN(n3347) );
  AOI22_X1 U3144 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[39] ), .B1(
        \dp/mul_feedback_exe_mem_int[40] ), .B2(n5186), .ZN(n3348) );
  NAND2_X1 U3145 ( .A1(n3347), .A2(n3348), .ZN(n6236) );
  AOI22_X1 U3146 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[47] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[47] ), .ZN(n3349) );
  AOI22_X1 U3147 ( .A1(n3943), .A2(\dp/a_neg_mult_id_exe_int[46] ), .B1(
        \dp/mul_feedback_exe_mem_int[47] ), .B2(n5186), .ZN(n3350) );
  NAND2_X1 U3148 ( .A1(n3349), .A2(n3350), .ZN(n6252) );
  AOI22_X1 U3149 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/a_shiftn[50] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[51] ), .ZN(n3351) );
  NAND2_X1 U3150 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[51] ), .A2(n3946), 
        .ZN(n3352) );
  OAI21_X1 U3151 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[51] ), .A(n3352), 
        .ZN(n3353) );
  AOI21_X1 U3152 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[50] ), 
        .A(n3353), .ZN(n3354) );
  NAND2_X1 U3153 ( .A1(n3351), .A2(n3354), .ZN(n6274) );
  NAND2_X1 U3154 ( .A1(n5145), .A2(n3900), .ZN(n3355) );
  NOR2_X1 U3155 ( .A1(n5685), .A2(n3355), .ZN(n5187) );
  INV_X1 U3156 ( .A(n5091), .ZN(n3356) );
  AOI21_X1 U3157 ( .B1(n5923), .B2(n5092), .A(n3356), .ZN(n3357) );
  XNOR2_X1 U3158 ( .A(n5925), .B(n5926), .ZN(n3358) );
  XNOR2_X1 U3159 ( .A(n3358), .B(n3357), .ZN(n3359) );
  INV_X1 U3160 ( .A(n3940), .ZN(n3360) );
  INV_X1 U3161 ( .A(n3923), .ZN(n3361) );
  AOI221_X1 U3162 ( .B1(n7069), .B2(n3923), .C1(n3360), .C2(n3361), .A(
        \intadd_1/B[11] ), .ZN(n3362) );
  NOR2_X1 U3163 ( .A1(\intadd_1/SUM[11] ), .A2(n7066), .ZN(n3363) );
  AOI211_X1 U3164 ( .C1(n3954), .C2(\dp/exs/alu_unit/shifter_out[12] ), .A(
        n3362), .B(n3363), .ZN(n3364) );
  INV_X1 U3165 ( .A(n6157), .ZN(n3365) );
  NAND3_X1 U3166 ( .A1(n3923), .A2(\intadd_1/B[11] ), .A3(n3365), .ZN(n3366)
         );
  OAI211_X1 U3167 ( .C1(n6027), .C2(n3359), .A(n3364), .B(n3366), .ZN(n6443)
         );
  NOR2_X1 U3168 ( .A1(n5230), .A2(n377), .ZN(n3367) );
  AOI21_X1 U3169 ( .B1(\dp/ids/rp1[19] ), .B2(n4136), .A(n3367), .ZN(n6826) );
  INV_X1 U3170 ( .A(n7056), .ZN(n3368) );
  NAND2_X1 U3171 ( .A1(\dp/a_mult_id_exe_int[13] ), .A2(n3876), .ZN(n3369) );
  OAI21_X1 U3172 ( .B1(n3368), .B2(n6847), .A(n3369), .ZN(n2933) );
  AOI22_X1 U3173 ( .A1(\dp/id_exe_regs/b_mult_reg/q[24] ), .A2(n3947), .B1(
        \dp/id_exe_regs/b_mult_reg/q[22] ), .B2(n3898), .ZN(n3370) );
  AOI22_X1 U3174 ( .A1(\dp/ids/rp2[23] ), .A2(n5213), .B1(rs_id[2]), .B2(n4648), .ZN(n3371) );
  NAND3_X1 U3175 ( .A1(n6958), .A2(n3370), .A3(n3371), .ZN(n2694) );
  INV_X1 U3176 ( .A(n4043), .ZN(n3372) );
  NAND2_X1 U3177 ( .A1(\dp/mul_feedback_exe_mem_int[31] ), .A2(n4016), .ZN(
        n3373) );
  OAI21_X1 U3178 ( .B1(n4043), .B2(\dp/b_adder_id_exe_int[31] ), .A(n4041), 
        .ZN(n3374) );
  NAND2_X1 U3179 ( .A1(n3374), .A2(n3373), .ZN(n3375) );
  OAI21_X1 U3180 ( .B1(wp_data[31]), .B2(n3372), .A(n3375), .ZN(n6161) );
  AOI22_X1 U3181 ( .A1(n5184), .A2(\dp/a_neg_mult_id_exe_int[46] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[46] ), .ZN(n3376) );
  AOI22_X1 U3182 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[45] ), .B1(
        \dp/mul_feedback_exe_mem_int[46] ), .B2(n5186), .ZN(n3377) );
  NAND2_X1 U3183 ( .A1(n3376), .A2(n3377), .ZN(n6250) );
  AOI22_X1 U3184 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/a_shiftn[48] ), .B1(
        n3946), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[49] ), .ZN(n3378) );
  NAND2_X1 U3185 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[49] ), .A2(n3945), .ZN(
        n3379) );
  OAI21_X1 U3186 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[49] ), .A(n3379), 
        .ZN(n3380) );
  AOI21_X1 U3187 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[48] ), 
        .A(n3380), .ZN(n3381) );
  NAND2_X1 U3188 ( .A1(n3378), .A2(n3381), .ZN(n6267) );
  AOI22_X1 U3189 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[56] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[56] ), .ZN(n3382) );
  AOI22_X1 U3190 ( .A1(n3943), .A2(\dp/a_neg_mult_id_exe_int[55] ), .B1(
        \dp/mul_feedback_exe_mem_int[56] ), .B2(n5186), .ZN(n3383) );
  NAND2_X1 U3191 ( .A1(n3382), .A2(n3383), .ZN(n6288) );
  AOI22_X1 U3192 ( .A1(n6326), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[58] ), 
        .B1(n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[59] ), .ZN(n3384) );
  NAND2_X1 U3193 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[59] ), .A2(n5188), 
        .ZN(n3385) );
  OAI21_X1 U3194 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[59] ), .A(n3385), 
        .ZN(n3386) );
  AOI21_X1 U3195 ( .B1(n5189), .B2(\dp/exs/alu_unit/mult/a_shiftn[58] ), .A(
        n3386), .ZN(n3387) );
  NAND2_X1 U3196 ( .A1(n3384), .A2(n3387), .ZN(n6295) );
  AOI22_X1 U3197 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[18] ), .A2(n3945), .B1(
        n5154), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[17] ), .ZN(n3388) );
  AOI22_X1 U3198 ( .A1(n3946), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[18] ), 
        .B1(n5189), .B2(\dp/exs/alu_unit/mult/a_shiftn[17] ), .ZN(n3389) );
  NAND2_X1 U3199 ( .A1(n6327), .A2(n4267), .ZN(n3390) );
  NAND3_X1 U3200 ( .A1(n3390), .A2(n3388), .A3(n3389), .ZN(n5970) );
  NAND2_X1 U3201 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[12] ), .A2(n6326), 
        .ZN(n3391) );
  AOI22_X1 U3202 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/a_shiftn[12] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[13] ), .ZN(n3392) );
  AOI21_X1 U3203 ( .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[13] ), .B2(n3946), 
        .A(n5688), .ZN(n3393) );
  NAND3_X1 U3204 ( .A1(n3391), .A2(n3392), .A3(n3393), .ZN(n5928) );
  AOI22_X1 U3205 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/ax2_shiftn[10] ), 
        .B1(n3945), .B2(\dp/exs/alu_unit/mult/ax2_shiftn[11] ), .ZN(n3394) );
  NAND2_X1 U3206 ( .A1(\dp/exs/alu_unit/mult/neg_ax2_shiftn[10] ), .A2(n6326), 
        .ZN(n3395) );
  OAI21_X1 U3207 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[10] ), .A(n3395), 
        .ZN(n3396) );
  AOI21_X1 U3208 ( .B1(n3946), .B2(\dp/exs/alu_unit/mult/neg_ax2_shiftn[11] ), 
        .A(n3396), .ZN(n3397) );
  NAND2_X1 U3209 ( .A1(n3394), .A2(n3397), .ZN(n5918) );
  AOI22_X1 U3210 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/ax2_shiftn[8] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/ax2_shiftn[9] ), .ZN(n3398) );
  NAND2_X1 U3211 ( .A1(\dp/exs/alu_unit/mult/neg_ax2_shiftn[8] ), .A2(n6326), 
        .ZN(n3399) );
  OAI21_X1 U3212 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[8] ), .A(n3399), .ZN(
        n3400) );
  AOI21_X1 U3213 ( .B1(n3946), .B2(\dp/exs/alu_unit/mult/neg_ax2_shiftn[9] ), 
        .A(n3400), .ZN(n3401) );
  NAND2_X1 U3214 ( .A1(n3398), .A2(n3401), .ZN(n5898) );
  XNOR2_X1 U3215 ( .A(n6098), .B(n6099), .ZN(n3402) );
  XNOR2_X1 U3216 ( .A(n3402), .B(n6100), .ZN(n3403) );
  INV_X1 U3217 ( .A(n6096), .ZN(n3404) );
  AOI221_X1 U3218 ( .B1(n7080), .B2(n6096), .C1(n7069), .C2(n3404), .A(
        \intadd_1/B[26] ), .ZN(n3405) );
  AOI21_X1 U3219 ( .B1(n3954), .B2(\dp/exs/alu_unit/shifter_out[27] ), .A(
        n3405), .ZN(n3406) );
  NAND3_X1 U3220 ( .A1(\intadd_1/B[26] ), .A2(n3952), .A3(n3404), .ZN(n3407)
         );
  OAI211_X1 U3221 ( .C1(\intadd_1/SUM[26] ), .C2(n7066), .A(n3406), .B(n3407), 
        .ZN(n3408) );
  AOI21_X1 U3222 ( .B1(n3403), .B2(n7076), .A(n3408), .ZN(n6417) );
  NOR2_X1 U3223 ( .A1(n5230), .A2(n367), .ZN(n3409) );
  AOI21_X1 U3224 ( .B1(\dp/ids/rp1[9] ), .B2(n4136), .A(n3409), .ZN(n6855) );
  INV_X1 U3225 ( .A(n5200), .ZN(n3410) );
  NAND2_X1 U3226 ( .A1(\dp/a_mult_id_exe_int[12] ), .A2(n3878), .ZN(n3411) );
  OAI21_X1 U3227 ( .B1(n3410), .B2(n6849), .A(n3411), .ZN(n2934) );
  AOI22_X1 U3228 ( .A1(\dp/id_exe_regs/b_mult_reg/q[21] ), .A2(n3956), .B1(
        \dp/id_exe_regs/b_mult_reg/q[19] ), .B2(n3896), .ZN(n3412) );
  AOI22_X1 U3229 ( .A1(rt_id[4]), .A2(n4648), .B1(\dp/ids/rp2[20] ), .B2(n5213), .ZN(n3413) );
  NAND3_X1 U3230 ( .A1(n3412), .A2(n6958), .A3(n3413), .ZN(n2697) );
  INV_X1 U3231 ( .A(\dp/mul_feedback_exe_mem_int[31] ), .ZN(n3414) );
  NAND2_X1 U3232 ( .A1(n5330), .A2(wp_data[31]), .ZN(n3415) );
  OAI21_X1 U3233 ( .B1(n3414), .B2(n5123), .A(n3415), .ZN(n7189) );
  AOI22_X1 U3234 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/a_shiftn[46] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[47] ), .ZN(n3416) );
  NAND2_X1 U3235 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[47] ), .A2(n3946), 
        .ZN(n3417) );
  OAI21_X1 U3236 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[47] ), .A(n3417), 
        .ZN(n3418) );
  AOI21_X1 U3237 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[46] ), 
        .A(n3418), .ZN(n3419) );
  NAND2_X1 U3238 ( .A1(n3416), .A2(n3419), .ZN(n6253) );
  AOI22_X1 U3239 ( .A1(n3946), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[53] ), 
        .B1(n6298), .B2(\dp/exs/alu_unit/mult/a_shiftn[52] ), .ZN(n3420) );
  NAND2_X1 U3240 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[52] ), .A2(n6326), 
        .ZN(n3421) );
  OAI21_X1 U3241 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[53] ), .A(n3421), 
        .ZN(n3422) );
  AOI21_X1 U3242 ( .B1(n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[53] ), .A(
        n3422), .ZN(n3423) );
  NAND2_X1 U3243 ( .A1(n3420), .A2(n3423), .ZN(n6279) );
  AOI22_X1 U3244 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[57] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[57] ), .ZN(n3424) );
  AOI22_X1 U3245 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[56] ), .B1(
        \dp/mul_feedback_exe_mem_int[57] ), .B2(n5156), .ZN(n3425) );
  NAND2_X1 U3246 ( .A1(n3424), .A2(n3425), .ZN(n6290) );
  AOI22_X1 U3247 ( .A1(n3943), .A2(\dp/a_neg_mult_id_exe_int[16] ), .B1(n5184), 
        .B2(\dp/a_neg_mult_id_exe_int[17] ), .ZN(n3426) );
  AOI22_X1 U3248 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[17] ), .B1(
        \dp/mul_feedback_exe_mem_int[17] ), .B2(n5186), .ZN(n3427) );
  NAND2_X1 U3249 ( .A1(n3426), .A2(n3427), .ZN(n5955) );
  AOI22_X1 U3250 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/ax2_shiftn[7] ), .B1(
        n5188), .B2(\dp/exs/alu_unit/mult/neg_ax2_shiftn[8] ), .ZN(n3428) );
  NAND2_X1 U3251 ( .A1(\dp/exs/alu_unit/mult/ax2_shiftn[8] ), .A2(n5187), .ZN(
        n3429) );
  OAI21_X1 U3252 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[7] ), .A(n3429), .ZN(
        n3430) );
  AOI21_X1 U3253 ( .B1(n5154), .B2(\dp/exs/alu_unit/mult/neg_ax2_shiftn[7] ), 
        .A(n3430), .ZN(n3431) );
  NAND2_X1 U3254 ( .A1(n3428), .A2(n3431), .ZN(n5886) );
  AOI21_X1 U3255 ( .B1(instr_if[31]), .B2(n3962), .A(n5637), .ZN(n3432) );
  NAND4_X1 U3256 ( .A1(n3929), .A2(n5602), .A3(n3432), .A4(n5614), .ZN(n3433)
         );
  NAND2_X1 U3257 ( .A1(n5652), .A2(n3433), .ZN(n5598) );
  INV_X1 U3258 ( .A(n6022), .ZN(n3434) );
  OAI21_X1 U3259 ( .B1(n5068), .B2(n3434), .A(n5067), .ZN(n3435) );
  XOR2_X1 U3260 ( .A(n6029), .B(n6030), .Z(n3436) );
  XNOR2_X1 U3261 ( .A(n3435), .B(n3436), .ZN(n3437) );
  NOR2_X1 U3262 ( .A1(n4730), .A2(n5243), .ZN(n3438) );
  NAND3_X1 U3263 ( .A1(\intadd_1/B[21] ), .A2(n3438), .A3(n3952), .ZN(n3439)
         );
  INV_X1 U3264 ( .A(n7080), .ZN(n3440) );
  AOI21_X1 U3265 ( .B1(n7069), .B2(n3438), .A(\intadd_1/B[21] ), .ZN(n3441) );
  OAI21_X1 U3266 ( .B1(n3438), .B2(n3440), .A(n3441), .ZN(n3442) );
  OAI211_X1 U3267 ( .C1(\intadd_1/SUM[21] ), .C2(n7066), .A(n3439), .B(n3442), 
        .ZN(n3443) );
  AOI21_X1 U3268 ( .B1(n7083), .B2(\dp/exs/alu_unit/shifter_out[22] ), .A(
        n3443), .ZN(n3444) );
  OAI21_X1 U3269 ( .B1(n6027), .B2(n3437), .A(n3444), .ZN(n6423) );
  NOR2_X1 U3270 ( .A1(n5230), .A2(n370), .ZN(n3445) );
  AOI21_X1 U3271 ( .B1(\dp/ids/rp1[12] ), .B2(n4136), .A(n3445), .ZN(n6849) );
  AND2_X1 U3272 ( .A1(\ctrl_u/curr_exe[0] ), .A2(n5667), .ZN(n3446) );
  OAI221_X1 U3273 ( .B1(n3446), .B2(n7340), .C1(n3446), .C2(
        \ctrl_u/curr_mem[0] ), .A(rst_mem_wb_regs), .ZN(\ctrl_u/n480 ) );
  INV_X1 U3274 ( .A(n5201), .ZN(n3447) );
  NAND2_X1 U3275 ( .A1(\dp/a_mult_id_exe_int[11] ), .A2(n3876), .ZN(n3448) );
  OAI21_X1 U3276 ( .B1(n3447), .B2(n6851), .A(n3448), .ZN(n2935) );
  AOI22_X1 U3277 ( .A1(n5213), .A2(\dp/ids/rp2[24] ), .B1(rs_id[3]), .B2(n4648), .ZN(n3449) );
  NAND3_X1 U3278 ( .A1(n6957), .A2(n6958), .A3(n3449), .ZN(n2693) );
  AOI222_X1 U3279 ( .A1(n5170), .A2(n4292), .B1(n4016), .B2(n4109), .C1(n5274), 
        .C2(n4043), .ZN(n3450) );
  INV_X1 U3280 ( .A(n3450), .ZN(n6124) );
  OAI22_X1 U3281 ( .A1(n5123), .A2(n4064), .B1(n5284), .B2(n3950), .ZN(n7197)
         );
  OAI21_X1 U3282 ( .B1(n5089), .B2(n5092), .A(n5925), .ZN(n3451) );
  INV_X1 U3283 ( .A(n3451), .ZN(n4001) );
  AOI22_X1 U3284 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/a_shiftn[33] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[34] ), .ZN(n3452) );
  NAND2_X1 U3285 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[34] ), .A2(n3946), 
        .ZN(n3453) );
  OAI21_X1 U3286 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[34] ), .A(n3453), 
        .ZN(n3454) );
  AOI21_X1 U3287 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[33] ), 
        .A(n3454), .ZN(n3455) );
  NAND2_X1 U3288 ( .A1(n3452), .A2(n3455), .ZN(n6200) );
  AOI22_X1 U3289 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[49] ), .B1(n3919), 
        .B2(\dp/a_neg_mult_id_exe_int[48] ), .ZN(n3456) );
  AOI22_X1 U3290 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[49] ), .B1(
        \dp/mul_feedback_exe_mem_int[49] ), .B2(n5186), .ZN(n3457) );
  NAND2_X1 U3291 ( .A1(n3456), .A2(n3457), .ZN(n6268) );
  AOI22_X1 U3292 ( .A1(n3946), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[55] ), 
        .B1(n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[55] ), .ZN(n3458) );
  NAND2_X1 U3293 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[54] ), .A2(n5189), .ZN(
        n3459) );
  OAI21_X1 U3294 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[55] ), .A(n3459), 
        .ZN(n3460) );
  AOI21_X1 U3295 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[54] ), 
        .A(n3460), .ZN(n3461) );
  NAND2_X1 U3296 ( .A1(n3458), .A2(n3461), .ZN(n6286) );
  AOI22_X1 U3297 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[58] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[58] ), .ZN(n3462) );
  AOI22_X1 U3298 ( .A1(n3943), .A2(\dp/a_neg_mult_id_exe_int[57] ), .B1(
        \dp/mul_feedback_exe_mem_int[58] ), .B2(n5186), .ZN(n3463) );
  NAND2_X1 U3299 ( .A1(n3462), .A2(n3463), .ZN(n6293) );
  INV_X1 U3300 ( .A(\intadd_1/n128 ), .ZN(n3464) );
  AOI21_X1 U3301 ( .B1(n4729), .B2(\intadd_1/n190 ), .A(n3464), .ZN(n3465) );
  OAI21_X1 U3302 ( .B1(n4038), .B2(\intadd_1/B[10] ), .A(\intadd_1/n123 ), 
        .ZN(n3466) );
  XOR2_X1 U3303 ( .A(n3465), .B(n3466), .Z(\intadd_1/SUM[10] ) );
  AOI22_X1 U3304 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[8] ), .B1(n5184), 
        .B2(\dp/a_neg_mult_id_exe_int[9] ), .ZN(n3467) );
  AOI22_X1 U3305 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[9] ), .B1(
        \dp/mul_feedback_exe_mem_int[9] ), .B2(n5186), .ZN(n3468) );
  NAND2_X1 U3306 ( .A1(n3467), .A2(n3468), .ZN(n5908) );
  NOR2_X1 U3307 ( .A1(n4303), .A2(n5342), .ZN(n3469) );
  OAI221_X1 U3308 ( .B1(n5675), .B2(n3469), .C1(n5675), .C2(n4300), .A(n5097), 
        .ZN(n5417) );
  AOI22_X1 U3309 ( .A1(n3931), .A2(\dp/ifs/pc_btb[19] ), .B1(
        btb_cache_read_address[19]), .B2(n5193), .ZN(n3470) );
  OAI21_X1 U3310 ( .B1(n3873), .B2(n4101), .A(n3470), .ZN(n6395) );
  NAND3_X1 U3311 ( .A1(\intadd_1/B[22] ), .A2(n3952), .A3(n6036), .ZN(n3471)
         );
  OAI21_X1 U3312 ( .B1(\intadd_1/B[22] ), .B2(n6037), .A(n3471), .ZN(n3472) );
  AOI21_X1 U3313 ( .B1(n4206), .B2(n6022), .A(n5032), .ZN(n3473) );
  XNOR2_X1 U3314 ( .A(n6040), .B(n6039), .ZN(n3474) );
  NAND2_X1 U3315 ( .A1(n3473), .A2(n3474), .ZN(n3475) );
  OAI211_X1 U3316 ( .C1(n3473), .C2(n3474), .A(n7076), .B(n3475), .ZN(n3476)
         );
  OAI21_X1 U3317 ( .B1(\intadd_1/SUM[22] ), .B2(n7066), .A(n3476), .ZN(n3477)
         );
  AOI211_X1 U3318 ( .C1(n3954), .C2(\dp/exs/alu_unit/shifter_out[23] ), .A(
        n3472), .B(n3477), .ZN(n6421) );
  XOR2_X1 U3319 ( .A(n5756), .B(n5757), .Z(n3478) );
  OAI21_X1 U3320 ( .B1(n5758), .B2(n3478), .A(n7076), .ZN(n3479) );
  AOI21_X1 U3321 ( .B1(n5758), .B2(n3478), .A(n3479), .ZN(n3480) );
  INV_X1 U3322 ( .A(n5752), .ZN(n3481) );
  NAND3_X1 U3323 ( .A1(\intadd_1/B[15] ), .A2(n3952), .A3(n3481), .ZN(n3482)
         );
  AOI221_X1 U3324 ( .B1(n7080), .B2(n5752), .C1(n7069), .C2(n3481), .A(
        \intadd_1/B[15] ), .ZN(n3483) );
  INV_X1 U3325 ( .A(n3483), .ZN(n3484) );
  OAI211_X1 U3326 ( .C1(\intadd_1/SUM[15] ), .C2(n7066), .A(n3482), .B(n3484), 
        .ZN(n3485) );
  AOI211_X1 U3327 ( .C1(n3954), .C2(\dp/exs/alu_unit/shifter_out[16] ), .A(
        n3480), .B(n3485), .ZN(n7437) );
  NOR2_X1 U3328 ( .A1(n5230), .A2(n366), .ZN(n3486) );
  AOI21_X1 U3329 ( .B1(\dp/ids/rp1[8] ), .B2(n4136), .A(n3486), .ZN(n6857) );
  AND2_X1 U3330 ( .A1(\ctrl_u/curr_exe[1] ), .A2(n5667), .ZN(n3487) );
  OAI221_X1 U3331 ( .B1(n3487), .B2(n7340), .C1(n3487), .C2(
        \ctrl_u/curr_mem[1] ), .A(rst_mem_wb_regs), .ZN(\ctrl_u/n479 ) );
  AOI21_X1 U3332 ( .B1(instr_if[3]), .B2(n5464), .A(n5463), .ZN(n3488) );
  OAI211_X1 U3333 ( .C1(n5594), .C2(n3488), .A(n5016), .B(n5474), .ZN(n3489)
         );
  OAI21_X1 U3334 ( .B1(n4485), .B2(n5599), .A(n3489), .ZN(n3490) );
  NAND2_X1 U3335 ( .A1(n3490), .A2(n3929), .ZN(\ctrl_u/n514 ) );
  INV_X1 U3336 ( .A(n5200), .ZN(n3491) );
  NAND2_X1 U3337 ( .A1(\dp/a_mult_id_exe_int[10] ), .A2(n3877), .ZN(n3492) );
  OAI21_X1 U3338 ( .B1(n3491), .B2(n6853), .A(n3492), .ZN(n2936) );
  NAND2_X1 U3339 ( .A1(n3947), .A2(n4388), .ZN(n3493) );
  OAI211_X1 U3340 ( .C1(n4820), .C2(n7047), .A(n6900), .B(n3493), .ZN(n2714)
         );
  NAND2_X1 U3341 ( .A1(n6991), .A2(rs_id[3]), .ZN(n3494) );
  AOI22_X1 U3342 ( .A1(\dp/b_adder_id_exe_int[24] ), .A2(n5210), .B1(
        \dp/ids/rp2[24] ), .B2(n3881), .ZN(n3495) );
  NAND3_X1 U3343 ( .A1(n3494), .A2(n3495), .A3(n6993), .ZN(n2661) );
  AOI222_X1 U3344 ( .A1(n5170), .A2(n4294), .B1(n4016), .B2(n4067), .C1(n5282), 
        .C2(n4024), .ZN(n3496) );
  INV_X1 U3345 ( .A(n3496), .ZN(n6105) );
  INV_X1 U3346 ( .A(n5006), .ZN(n3497) );
  AOI22_X1 U3347 ( .A1(n6004), .A2(n6005), .B1(n4904), .B2(n3497), .ZN(n4902)
         );
  OAI22_X1 U3348 ( .A1(n3950), .A2(n5301), .B1(n4081), .B2(n5123), .ZN(n7221)
         );
  OAI22_X1 U3349 ( .A1(n5172), .A2(n5310), .B1(n4074), .B2(n5173), .ZN(n7231)
         );
  AOI22_X1 U3350 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[59] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[59] ), .ZN(n3498) );
  AOI22_X1 U3351 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[58] ), .B1(
        \dp/mul_feedback_exe_mem_int[59] ), .B2(n5156), .ZN(n3499) );
  NAND2_X1 U3352 ( .A1(n3498), .A2(n3499), .ZN(n6296) );
  NAND2_X1 U3353 ( .A1(n6147), .A2(n6148), .ZN(n3500) );
  OAI21_X1 U3354 ( .B1(n3500), .B2(n6308), .A(n4869), .ZN(n6311) );
  AOI22_X1 U3355 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/a_shiftn[61] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[62] ), .ZN(n3501) );
  NAND2_X1 U3356 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[62] ), .A2(n3946), 
        .ZN(n3502) );
  OAI21_X1 U3357 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[62] ), .A(n3502), 
        .ZN(n3503) );
  AOI21_X1 U3358 ( .B1(n5154), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[61] ), 
        .A(n3503), .ZN(n3504) );
  NAND2_X1 U3359 ( .A1(n3501), .A2(n3504), .ZN(n6305) );
  AOI22_X1 U3360 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[13] ), .B1(n5184), 
        .B2(\dp/a_neg_mult_id_exe_int[14] ), .ZN(n3505) );
  AOI22_X1 U3361 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[14] ), .B1(
        \dp/mul_feedback_exe_mem_int[14] ), .B2(n5186), .ZN(n3506) );
  NAND2_X1 U3362 ( .A1(n3505), .A2(n3506), .ZN(n5939) );
  AOI22_X1 U3363 ( .A1(n5188), .A2(\dp/exs/alu_unit/mult/neg_ax2_shiftn[7] ), 
        .B1(n5187), .B2(\dp/exs/alu_unit/mult/ax2_shiftn[7] ), .ZN(n3507) );
  NAND3_X1 U3364 ( .A1(n5690), .A2(n5691), .A3(n3507), .ZN(n5874) );
  INV_X1 U3365 ( .A(n4052), .ZN(n3508) );
  NAND3_X1 U3366 ( .A1(n4933), .A2(n5480), .A3(n3508), .ZN(n5547) );
  AOI22_X1 U3367 ( .A1(\dp/ifs/pc_btb[20] ), .A2(n3931), .B1(
        btb_cache_read_address[20]), .B2(n5193), .ZN(n3509) );
  INV_X1 U3368 ( .A(n3509), .ZN(n4877) );
  INV_X1 U3369 ( .A(n5109), .ZN(n3510) );
  AOI221_X1 U3370 ( .B1(n7069), .B2(n5109), .C1(n7080), .C2(n3510), .A(
        \intadd_1/B[10] ), .ZN(n3511) );
  XOR2_X1 U3371 ( .A(n5923), .B(n5921), .Z(n3512) );
  NAND2_X1 U3372 ( .A1(n5922), .A2(n3512), .ZN(n3513) );
  OAI211_X1 U3373 ( .C1(n5922), .C2(n3512), .A(n7076), .B(n3513), .ZN(n3514)
         );
  NAND3_X1 U3374 ( .A1(\intadd_1/B[10] ), .A2(n5109), .A3(n3952), .ZN(n3515)
         );
  OAI211_X1 U3375 ( .C1(\intadd_1/SUM[10] ), .C2(n7066), .A(n3514), .B(n3515), 
        .ZN(n3516) );
  AOI211_X1 U3376 ( .C1(n7083), .C2(\dp/exs/alu_unit/shifter_out[11] ), .A(
        n3511), .B(n3516), .ZN(n6445) );
  NOR2_X1 U3377 ( .A1(n5230), .A2(n368), .ZN(n3517) );
  AOI21_X1 U3378 ( .B1(\dp/ids/rp1[10] ), .B2(n4136), .A(n3517), .ZN(n6853) );
  AND2_X1 U3379 ( .A1(\ctrl_u/curr_exe[5] ), .A2(n5667), .ZN(n3518) );
  OAI221_X1 U3380 ( .B1(n3518), .B2(n7340), .C1(n3518), .C2(
        \ctrl_u/curr_mem[5] ), .A(rst_mem_wb_regs), .ZN(\ctrl_u/n475 ) );
  OAI21_X1 U3381 ( .B1(\ctrl_u/n66 ), .B2(n5599), .A(n5598), .ZN(\ctrl_u/n518 ) );
  INV_X1 U3382 ( .A(n5201), .ZN(n3519) );
  NAND2_X1 U3383 ( .A1(\dp/a_mult_id_exe_int[9] ), .A2(n3878), .ZN(n3520) );
  OAI21_X1 U3384 ( .B1(n3519), .B2(n6855), .A(n3520), .ZN(n2937) );
  AOI22_X1 U3385 ( .A1(\dp/ids/rp2[5] ), .A2(n5213), .B1(\dp/imm_id_int[5] ), 
        .B2(n4675), .ZN(n3521) );
  AOI22_X1 U3386 ( .A1(n4142), .A2(n3947), .B1(n4388), .B2(n3896), .ZN(n3522)
         );
  NAND2_X1 U3387 ( .A1(n3521), .A2(n3522), .ZN(n2712) );
  NAND2_X1 U3388 ( .A1(n6991), .A2(rs_id[2]), .ZN(n3523) );
  AOI22_X1 U3389 ( .A1(\dp/b_adder_id_exe_int[23] ), .A2(n5209), .B1(
        \dp/ids/rp2[23] ), .B2(n3881), .ZN(n3524) );
  NAND3_X1 U3390 ( .A1(n3523), .A2(n3524), .A3(n6993), .ZN(n2662) );
  OAI22_X1 U3391 ( .A1(n5173), .A2(n4067), .B1(n5282), .B2(n5172), .ZN(n7195)
         );
  OAI22_X1 U3392 ( .A1(n4040), .A2(wp_data[7]), .B1(
        \dp/mul_feedback_exe_mem_int[7] ), .B2(n3922), .ZN(n3525) );
  AOI21_X1 U3393 ( .B1(n4341), .B2(n5135), .A(n3525), .ZN(n5882) );
  AOI22_X1 U3394 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[37] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[37] ), .ZN(n3526) );
  AOI22_X1 U3395 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[36] ), .B1(
        \dp/mul_feedback_exe_mem_int[37] ), .B2(n5186), .ZN(n3527) );
  NAND2_X1 U3396 ( .A1(n3526), .A2(n3527), .ZN(n6212) );
  AOI22_X1 U3397 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[41] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[41] ), .ZN(n3528) );
  AOI22_X1 U3398 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[40] ), .B1(
        \dp/mul_feedback_exe_mem_int[41] ), .B2(n5186), .ZN(n3529) );
  NAND2_X1 U3399 ( .A1(n3528), .A2(n3529), .ZN(n6239) );
  AOI22_X1 U3400 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/a_shiftn[41] ), .B1(
        n3946), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[42] ), .ZN(n3530) );
  NAND2_X1 U3401 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[41] ), .A2(n6326), 
        .ZN(n3531) );
  OAI21_X1 U3402 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[42] ), .A(n3531), 
        .ZN(n3532) );
  AOI21_X1 U3403 ( .B1(n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[42] ), .A(
        n3532), .ZN(n3533) );
  NAND2_X1 U3404 ( .A1(n3530), .A2(n3533), .ZN(n6243) );
  AOI22_X1 U3405 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/a_shiftn[47] ), .B1(
        n3946), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[48] ), .ZN(n3534) );
  NAND2_X1 U3406 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[48] ), .A2(n3945), .ZN(
        n3535) );
  OAI21_X1 U3407 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[48] ), .A(n3535), 
        .ZN(n3536) );
  AOI21_X1 U3408 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[47] ), 
        .A(n3536), .ZN(n3537) );
  NAND2_X1 U3409 ( .A1(n3534), .A2(n3537), .ZN(n6266) );
  AOI22_X1 U3410 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[51] ), .B1(n3919), 
        .B2(\dp/a_neg_mult_id_exe_int[50] ), .ZN(n3538) );
  AOI22_X1 U3411 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[51] ), .B1(
        \dp/mul_feedback_exe_mem_int[51] ), .B2(n5186), .ZN(n3539) );
  NAND2_X1 U3412 ( .A1(n3538), .A2(n3539), .ZN(n6273) );
  AOI22_X1 U3413 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[60] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[60] ), .ZN(n3540) );
  AOI22_X1 U3414 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[59] ), .B1(
        \dp/mul_feedback_exe_mem_int[60] ), .B2(n5186), .ZN(n3541) );
  NAND2_X1 U3415 ( .A1(n3540), .A2(n3541), .ZN(n6299) );
  AOI22_X1 U3416 ( .A1(n3946), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[61] ), 
        .B1(n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[61] ), .ZN(n3542) );
  NAND2_X1 U3417 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[60] ), .A2(n6298), .ZN(
        n3543) );
  OAI21_X1 U3418 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[61] ), .A(n3543), 
        .ZN(n3544) );
  AOI21_X1 U3419 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[60] ), 
        .A(n3544), .ZN(n3545) );
  NAND2_X1 U3420 ( .A1(n3542), .A2(n3545), .ZN(n6302) );
  OAI211_X1 U3421 ( .C1(n5627), .C2(n5588), .A(n4844), .B(n4850), .ZN(n5549)
         );
  AOI22_X1 U3422 ( .A1(n4122), .A2(n4822), .B1(n4221), .B2(n4356), .ZN(n4746)
         );
  OAI21_X1 U3423 ( .B1(n6136), .B2(n4023), .A(n6135), .ZN(n3546) );
  OAI21_X1 U3424 ( .B1(n3547), .B2(n3548), .A(n3546), .ZN(n6119) );
  INV_X1 U3425 ( .A(n6148), .ZN(n3547) );
  INV_X1 U3426 ( .A(n6136), .ZN(n3548) );
  OR2_X1 U3427 ( .A1(n5922), .A2(n5921), .ZN(n5092) );
  AOI21_X1 U3428 ( .B1(\dp/exs/alu_unit/mult/ax2_shiftn[6] ), .B2(n5187), .A(
        n5692), .ZN(n3549) );
  AOI22_X1 U3429 ( .A1(\dp/exs/alu_unit/mult/neg_ax2_shiftn[6] ), .A2(n5188), 
        .B1(n6298), .B2(\dp/exs/alu_unit/mult/ax2_shiftn[5] ), .ZN(n3550) );
  NAND3_X1 U3430 ( .A1(n3549), .A2(n5693), .A3(n3550), .ZN(n5868) );
  OR2_X1 U3431 ( .A1(n6292), .A2(n6293), .ZN(n6685) );
  AOI22_X1 U3432 ( .A1(\dp/a_neg_mult_id_exe_int[2] ), .A2(n5184), .B1(
        \dp/mul_feedback_exe_mem_int[2] ), .B2(n5156), .ZN(n3551) );
  NAND3_X1 U3433 ( .A1(n5718), .A2(n6466), .A3(n3551), .ZN(n5814) );
  NOR4_X1 U3434 ( .A1(n5155), .A2(n5162), .A3(n5164), .A4(n5149), .ZN(n3552)
         );
  NAND3_X1 U3435 ( .A1(n5158), .A2(n7298), .A3(\ctrl_u/curr_exe[18] ), .ZN(
        n3553) );
  OAI211_X1 U3436 ( .C1(n3552), .C2(n4025), .A(n5753), .B(n3553), .ZN(n5755)
         );
  AOI21_X1 U3437 ( .B1(n5670), .B2(\ctrl_u/curr_mem[4] ), .A(n5229), .ZN(n7428) );
  INV_X1 U3438 ( .A(n3953), .ZN(n3554) );
  INV_X1 U3439 ( .A(n3992), .ZN(n3555) );
  AOI221_X1 U3440 ( .B1(n7080), .B2(n3992), .C1(n3554), .C2(n3555), .A(
        \intadd_1/B[9] ), .ZN(n3556) );
  XOR2_X1 U3441 ( .A(n5918), .B(n5917), .Z(n3557) );
  NAND2_X1 U3442 ( .A1(n3908), .A2(n3557), .ZN(n3558) );
  OAI211_X1 U3443 ( .C1(n3908), .C2(n3557), .A(n7076), .B(n3558), .ZN(n3559)
         );
  NAND3_X1 U3444 ( .A1(\intadd_1/B[9] ), .A2(n3952), .A3(n3555), .ZN(n3560) );
  OAI211_X1 U3445 ( .C1(\intadd_1/SUM[9] ), .C2(n7066), .A(n3559), .B(n3560), 
        .ZN(n3561) );
  AOI211_X1 U3446 ( .C1(\dp/exs/alu_unit/shifter_out[10] ), .C2(n3954), .A(
        n3556), .B(n3561), .ZN(n6447) );
  NOR2_X1 U3447 ( .A1(n5230), .A2(n363), .ZN(n3562) );
  AOI21_X1 U3448 ( .B1(\dp/ids/rp1[5] ), .B2(n4136), .A(n3562), .ZN(n6873) );
  INV_X1 U3449 ( .A(n5417), .ZN(n3563) );
  OAI21_X1 U3450 ( .B1(n5658), .B2(n3563), .A(n5674), .ZN(pc_en) );
  AOI211_X1 U3451 ( .C1(\dp/pc_plus4_out_if_int[25] ), .C2(n3936), .A(n6401), 
        .B(n5004), .ZN(n3564) );
  AOI21_X1 U3452 ( .B1(\dp/ifs/pc_btb[25] ), .B2(n3931), .A(n5047), .ZN(n3565)
         );
  NAND2_X1 U3453 ( .A1(n4901), .A2(n3884), .ZN(n3566) );
  NAND3_X1 U3454 ( .A1(n3566), .A2(n3564), .A3(n3565), .ZN(n2532) );
  AND2_X1 U3455 ( .A1(\ctrl_u/curr_exe[9] ), .A2(n5667), .ZN(n3567) );
  OAI221_X1 U3456 ( .B1(n3567), .B2(n7340), .C1(n3567), .C2(ld_type_mem[1]), 
        .A(rst_mem_wb_regs), .ZN(\ctrl_u/n471 ) );
  OAI21_X1 U3457 ( .B1(n4454), .B2(n5599), .A(n5598), .ZN(\ctrl_u/n543 ) );
  INV_X1 U3458 ( .A(n5202), .ZN(n3568) );
  NAND2_X1 U3459 ( .A1(\dp/a_mult_id_exe_int[8] ), .A2(n3877), .ZN(n3569) );
  OAI21_X1 U3460 ( .B1(n3568), .B2(n6857), .A(n3569), .ZN(n2938) );
  NAND2_X1 U3461 ( .A1(\dp/id_exe_regs/b_mult_reg/q[26] ), .A2(n3947), .ZN(
        n3570) );
  NAND2_X1 U3462 ( .A1(\dp/id_exe_regs/b_mult_reg/q[24] ), .A2(n3897), .ZN(
        n3571) );
  OAI211_X1 U3463 ( .C1(n6979), .C2(n4820), .A(n3570), .B(n3571), .ZN(n2692)
         );
  AOI22_X1 U3464 ( .A1(\dp/b_adder_id_exe_int[22] ), .A2(n5210), .B1(
        \dp/ids/rp2[22] ), .B2(n3880), .ZN(n3572) );
  NAND2_X1 U3465 ( .A1(n6991), .A2(rs_id[1]), .ZN(n3573) );
  NAND3_X1 U3466 ( .A1(n3573), .A2(n3572), .A3(n6993), .ZN(n2663) );
  OAI21_X1 U3467 ( .B1(n6134), .B2(n3574), .A(n3575), .ZN(n6137) );
  INV_X1 U3468 ( .A(n6141), .ZN(n3574) );
  INV_X1 U3469 ( .A(n6142), .ZN(n3575) );
  NOR2_X1 U3470 ( .A1(n4730), .A2(n5243), .ZN(n3576) );
  XOR2_X1 U3471 ( .A(n4225), .B(n3576), .Z(\intadd_1/A[21] ) );
  AOI22_X1 U3472 ( .A1(n5070), .A2(n5049), .B1(n4287), .B2(n5332), .ZN(n3577)
         );
  INV_X1 U3473 ( .A(n3577), .ZN(n4986) );
  OAI22_X1 U3474 ( .A1(n5173), .A2(n4089), .B1(n5299), .B2(n5172), .ZN(n7219)
         );
  OR2_X1 U3475 ( .A1(n5943), .A2(n5942), .ZN(n4814) );
  NAND2_X1 U3476 ( .A1(wp_data[9]), .A2(n5330), .ZN(n3578) );
  OAI21_X1 U3477 ( .B1(n4082), .B2(n5123), .A(n3578), .ZN(n7233) );
  AOI22_X1 U3478 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[32] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[32] ), .ZN(n3579) );
  AOI22_X1 U3479 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[31] ), .B1(
        \dp/mul_feedback_exe_mem_int[32] ), .B2(n5186), .ZN(n3580) );
  NAND2_X1 U3480 ( .A1(n3579), .A2(n3580), .ZN(n6312) );
  AOI22_X1 U3481 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[34] ), .B1(n3919), 
        .B2(\dp/a_neg_mult_id_exe_int[33] ), .ZN(n3581) );
  AOI22_X1 U3482 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[34] ), .B1(
        \dp/mul_feedback_exe_mem_int[34] ), .B2(n5186), .ZN(n3582) );
  NAND2_X1 U3483 ( .A1(n3581), .A2(n3582), .ZN(n6199) );
  AOI22_X1 U3484 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[36] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[36] ), .ZN(n3583) );
  AOI22_X1 U3485 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[35] ), .B1(
        \dp/mul_feedback_exe_mem_int[36] ), .B2(n5186), .ZN(n3584) );
  NAND2_X1 U3486 ( .A1(n3583), .A2(n3584), .ZN(n6210) );
  AOI22_X1 U3487 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[38] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[38] ), .ZN(n3585) );
  AOI22_X1 U3488 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[37] ), .B1(
        \dp/mul_feedback_exe_mem_int[38] ), .B2(n5186), .ZN(n3586) );
  NAND2_X1 U3489 ( .A1(n3585), .A2(n3586), .ZN(n6215) );
  AOI22_X1 U3490 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/a_shiftn[39] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[40] ), .ZN(n3587) );
  NAND2_X1 U3491 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[40] ), .A2(n3946), 
        .ZN(n3588) );
  OAI21_X1 U3492 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[40] ), .A(n3588), 
        .ZN(n3589) );
  AOI21_X1 U3493 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[39] ), 
        .A(n3589), .ZN(n3590) );
  NAND2_X1 U3494 ( .A1(n3587), .A2(n3590), .ZN(n6237) );
  AOI22_X1 U3495 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[41] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[42] ), .ZN(n3591) );
  AOI22_X1 U3496 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[42] ), .B1(
        \dp/mul_feedback_exe_mem_int[42] ), .B2(n5186), .ZN(n3592) );
  NAND2_X1 U3497 ( .A1(n3591), .A2(n3592), .ZN(n6242) );
  AOI22_X1 U3498 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[44] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[44] ), .ZN(n3593) );
  AOI22_X1 U3499 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[43] ), .B1(
        \dp/mul_feedback_exe_mem_int[44] ), .B2(n5186), .ZN(n3594) );
  NAND2_X1 U3500 ( .A1(n3593), .A2(n3594), .ZN(n6246) );
  AOI22_X1 U3501 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/a_shiftn[45] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[46] ), .ZN(n3595) );
  NAND2_X1 U3502 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[46] ), .A2(n3946), 
        .ZN(n3596) );
  OAI21_X1 U3503 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[46] ), .A(n3596), 
        .ZN(n3597) );
  AOI21_X1 U3504 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[45] ), 
        .A(n3597), .ZN(n3598) );
  NAND2_X1 U3505 ( .A1(n3595), .A2(n3598), .ZN(n6251) );
  AOI22_X1 U3506 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[48] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[48] ), .ZN(n3599) );
  AOI22_X1 U3507 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[47] ), .B1(
        \dp/mul_feedback_exe_mem_int[48] ), .B2(n5186), .ZN(n3600) );
  NAND2_X1 U3508 ( .A1(n3599), .A2(n3600), .ZN(n6265) );
  AOI22_X1 U3509 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[49] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[50] ), .ZN(n3601) );
  AOI22_X1 U3510 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[50] ), .B1(
        \dp/mul_feedback_exe_mem_int[50] ), .B2(n5186), .ZN(n3602) );
  NAND2_X1 U3511 ( .A1(n3601), .A2(n3602), .ZN(n6271) );
  AOI22_X1 U3512 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[52] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[52] ), .ZN(n3603) );
  AOI22_X1 U3513 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[51] ), .B1(
        \dp/mul_feedback_exe_mem_int[52] ), .B2(n5186), .ZN(n3604) );
  NAND2_X1 U3514 ( .A1(n3603), .A2(n3604), .ZN(n6276) );
  AOI22_X1 U3515 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[54] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[54] ), .ZN(n3605) );
  AOI22_X1 U3516 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[53] ), .B1(
        \dp/mul_feedback_exe_mem_int[54] ), .B2(n5186), .ZN(n3606) );
  NAND2_X1 U3517 ( .A1(n3605), .A2(n3606), .ZN(n6283) );
  AOI22_X1 U3518 ( .A1(n3946), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[58] ), 
        .B1(n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[58] ), .ZN(n3607) );
  NAND2_X1 U3519 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[57] ), .A2(n6326), 
        .ZN(n3608) );
  OAI21_X1 U3520 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[58] ), .A(n3608), 
        .ZN(n3609) );
  AOI21_X1 U3521 ( .B1(n6298), .B2(\dp/exs/alu_unit/mult/a_shiftn[57] ), .A(
        n3609), .ZN(n3610) );
  NAND2_X1 U3522 ( .A1(n3607), .A2(n3610), .ZN(n6292) );
  AOI22_X1 U3523 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[61] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[61] ), .ZN(n3611) );
  AOI22_X1 U3524 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[60] ), .B1(
        \dp/mul_feedback_exe_mem_int[61] ), .B2(n5186), .ZN(n3612) );
  NAND2_X1 U3525 ( .A1(n3611), .A2(n3612), .ZN(n6301) );
  INV_X1 U3526 ( .A(n5337), .ZN(n3613) );
  NOR2_X1 U3527 ( .A1(n5336), .A2(n3613), .ZN(n5822) );
  AOI222_X1 U3528 ( .A1(n5170), .A2(n4293), .B1(n4016), .B2(n4068), .C1(n5278), 
        .C2(n4043), .ZN(n3614) );
  INV_X1 U3529 ( .A(n3614), .ZN(n6113) );
  AOI21_X1 U3530 ( .B1(\intadd_1/n37 ), .B2(\intadd_1/n39 ), .A(\intadd_1/n36 ), .ZN(n3615) );
  NAND2_X1 U3531 ( .A1(\intadd_1/n33 ), .A2(n4229), .ZN(n3616) );
  XOR2_X1 U3532 ( .A(n3615), .B(n3616), .Z(\intadd_1/SUM[25] ) );
  AOI22_X1 U3533 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[9] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[10] ), .ZN(n3617) );
  AOI22_X1 U3534 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[10] ), .B1(
        \dp/mul_feedback_exe_mem_int[10] ), .B2(n5186), .ZN(n3618) );
  NAND2_X1 U3535 ( .A1(n3617), .A2(n3618), .ZN(n5917) );
  AOI22_X1 U3536 ( .A1(n6323), .A2(\dp/a_neg_mult_id_exe_int[5] ), .B1(n5184), 
        .B2(\dp/a_neg_mult_id_exe_int[6] ), .ZN(n3619) );
  AOI22_X1 U3537 ( .A1(n6322), .A2(\dp/a_mult_id_exe_int[6] ), .B1(
        \dp/mul_feedback_exe_mem_int[6] ), .B2(n5156), .ZN(n3620) );
  NAND2_X1 U3538 ( .A1(n3619), .A2(n3620), .ZN(n5152) );
  OR2_X1 U3539 ( .A1(n6295), .A2(n6296), .ZN(n6691) );
  NAND2_X1 U3540 ( .A1(n5352), .A2(rst_mem_wb_regs), .ZN(n3621) );
  OAI21_X1 U3541 ( .B1(n4821), .B2(n4876), .A(n3621), .ZN(n5349) );
  NAND3_X1 U3542 ( .A1(n4933), .A2(n4850), .A3(n5550), .ZN(n5557) );
  NOR2_X1 U3543 ( .A1(n4733), .A2(n3622), .ZN(n3623) );
  INV_X1 U3544 ( .A(n3623), .ZN(n3624) );
  AOI221_X1 U3545 ( .B1(n7080), .B2(n3623), .C1(n7069), .C2(n3624), .A(
        \intadd_1/B[0] ), .ZN(n3625) );
  AND3_X1 U3546 ( .A1(\intadd_1/B[0] ), .A2(n3952), .A3(n3624), .ZN(n3626) );
  AOI211_X1 U3547 ( .C1(\dp/exs/alu_unit/shifter_out[1] ), .C2(n3954), .A(
        n3625), .B(n3626), .ZN(n3627) );
  OAI211_X1 U3548 ( .C1(n6467), .C2(n6468), .A(n6466), .B(n7076), .ZN(n3628)
         );
  OAI211_X1 U3549 ( .C1(\intadd_1/SUM[0] ), .C2(n7066), .A(n3627), .B(n3628), 
        .ZN(n6470) );
  INV_X1 U3550 ( .A(n4715), .ZN(n3622) );
  NOR2_X1 U3551 ( .A1(n5230), .A2(n360), .ZN(n3629) );
  AOI21_X1 U3552 ( .B1(\dp/ids/rp1[2] ), .B2(n4136), .A(n3629), .ZN(n6884) );
  INV_X1 U3553 ( .A(\dp/ids/rp2[4] ), .ZN(n7045) );
  AND2_X1 U3554 ( .A1(\ctrl_u/curr_exe[11] ), .A2(n5667), .ZN(n3630) );
  OAI221_X1 U3555 ( .B1(n3630), .B2(n7340), .C1(n3630), .C2(
        \ctrl_u/curr_mem_11 ), .A(rst_mem_wb_regs), .ZN(\ctrl_u/n469 ) );
  OAI21_X1 U3556 ( .B1(\ctrl_u/n72 ), .B2(n5599), .A(n5598), .ZN(\ctrl_u/n550 ) );
  NOR2_X1 U3557 ( .A1(n4028), .A2(n5009), .ZN(n3631) );
  OAI211_X1 U3558 ( .C1(n3937), .C2(n5087), .A(n4004), .B(n3631), .ZN(n3041)
         );
  AOI22_X1 U3559 ( .A1(n3883), .A2(n4900), .B1(n3895), .B2(\dp/ifs/pc_btb[21] ), .ZN(n3632) );
  AOI211_X1 U3560 ( .C1(n7108), .C2(btb_cache_read_address[21]), .A(n6400), 
        .B(n4311), .ZN(n3633) );
  NAND2_X1 U3561 ( .A1(n3632), .A2(n3633), .ZN(n2536) );
  INV_X1 U3562 ( .A(n5201), .ZN(n3634) );
  NAND2_X1 U3563 ( .A1(\dp/a_mult_id_exe_int[3] ), .A2(n3877), .ZN(n3635) );
  OAI21_X1 U3564 ( .B1(n3634), .B2(n6882), .A(n3635), .ZN(n2943) );
  NAND2_X1 U3565 ( .A1(n5147), .A2(n3896), .ZN(n3636) );
  NAND2_X1 U3566 ( .A1(n4393), .A2(n5211), .ZN(n3637) );
  OAI211_X1 U3567 ( .C1(n7052), .C2(n4820), .A(n3636), .B(n3637), .ZN(n2715)
         );
  NAND2_X1 U3568 ( .A1(\dp/ids/rp2[21] ), .A2(n3880), .ZN(n3638) );
  NAND2_X1 U3569 ( .A1(\dp/b_adder_id_exe_int[21] ), .A2(n5206), .ZN(n3639) );
  NAND4_X1 U3570 ( .A1(n6993), .A2(n6985), .A3(n3638), .A4(n3639), .ZN(n2664)
         );
  INV_X1 U3571 ( .A(n5106), .ZN(n3640) );
  AOI22_X1 U3572 ( .A1(n4106), .A2(n5101), .B1(n5104), .B2(n3640), .ZN(n3641)
         );
  NAND2_X1 U3574 ( .A1(\intadd_1/n70 ), .A2(n5060), .ZN(n3643) );
  OAI211_X1 U3575 ( .C1(\intadd_1/n69 ), .C2(\intadd_1/n89 ), .A(n5059), .B(
        n3643), .ZN(n5058) );
  OAI22_X1 U3576 ( .A1(n5173), .A2(n4063), .B1(n5314), .B2(n5171), .ZN(n7235)
         );
  AOI22_X1 U3577 ( .A1(n6326), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[36] ), 
        .B1(n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[37] ), .ZN(n3644) );
  NAND2_X1 U3578 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[37] ), .A2(n3946), 
        .ZN(n3645) );
  OAI21_X1 U3579 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[37] ), .A(n3645), 
        .ZN(n3646) );
  AOI21_X1 U3580 ( .B1(n5189), .B2(\dp/exs/alu_unit/mult/a_shiftn[36] ), .A(
        n3646), .ZN(n3647) );
  NAND2_X1 U3581 ( .A1(n3644), .A2(n3647), .ZN(n6213) );
  AOI22_X1 U3582 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/a_shiftn[38] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[39] ), .ZN(n3648) );
  NAND2_X1 U3583 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[39] ), .A2(n3946), 
        .ZN(n3649) );
  OAI21_X1 U3584 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[39] ), .A(n3649), 
        .ZN(n3650) );
  AOI21_X1 U3585 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[38] ), 
        .A(n3650), .ZN(n3651) );
  NAND2_X1 U3586 ( .A1(n3648), .A2(n3651), .ZN(n6217) );
  INV_X1 U3587 ( .A(n6542), .ZN(n3652) );
  AOI21_X1 U3588 ( .B1(n6554), .B2(n6551), .A(n6555), .ZN(n3653) );
  OAI21_X1 U3589 ( .B1(n6241), .B2(n3652), .A(n3653), .ZN(n6561) );
  INV_X1 U3590 ( .A(n6605), .ZN(n3654) );
  AOI21_X1 U3591 ( .B1(n6616), .B2(n6613), .A(n6617), .ZN(n3655) );
  OAI21_X1 U3592 ( .B1(n6270), .B2(n3654), .A(n3655), .ZN(n6623) );
  AOI22_X1 U3593 ( .A1(n4776), .A2(n4709), .B1(\intadd_1/B[26] ), .B2(
        \intadd_1/A[26] ), .ZN(n4775) );
  AOI22_X1 U3594 ( .A1(n5041), .A2(n5040), .B1(\intadd_2/A[4] ), .B2(n4210), 
        .ZN(n5039) );
  NOR2_X1 U3595 ( .A1(taken), .A2(btb_cache_data_out_rw[31]), .ZN(n3656) );
  NOR2_X1 U3596 ( .A1(n6168), .A2(n3656), .ZN(n6169) );
  AOI22_X1 U3597 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/a_shiftn[28] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[29] ), .ZN(n3657) );
  NAND2_X1 U3598 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[29] ), .A2(n5188), 
        .ZN(n3658) );
  OAI21_X1 U3599 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[29] ), .A(n3658), 
        .ZN(n3659) );
  AOI21_X1 U3600 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[28] ), 
        .A(n3659), .ZN(n3660) );
  NAND2_X1 U3601 ( .A1(n3657), .A2(n3660), .ZN(n6141) );
  INV_X1 U3602 ( .A(\intadd_1/B[25] ), .ZN(n3661) );
  INV_X1 U3603 ( .A(n6082), .ZN(n3662) );
  OAI221_X1 U3604 ( .B1(n6082), .B2(n7080), .C1(n3662), .C2(n7069), .A(n3661), 
        .ZN(n3663) );
  OAI221_X1 U3605 ( .B1(n3661), .B2(n6082), .C1(n3661), .C2(n3952), .A(n3663), 
        .ZN(n6083) );
  AOI222_X1 U3606 ( .A1(n3903), .A2(n4308), .B1(n5136), .B2(n4089), .C1(n4024), 
        .C2(n5299), .ZN(n3664) );
  INV_X1 U3607 ( .A(n3664), .ZN(n5752) );
  INV_X1 U3608 ( .A(n5931), .ZN(n3665) );
  OAI21_X1 U3609 ( .B1(n4950), .B2(n3665), .A(n4951), .ZN(n5945) );
  AOI22_X1 U3610 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[11] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[12] ), .ZN(n3666) );
  AOI22_X1 U3611 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[12] ), .B1(
        \dp/mul_feedback_exe_mem_int[12] ), .B2(n5186), .ZN(n3667) );
  NAND2_X1 U3612 ( .A1(n3666), .A2(n3667), .ZN(n5926) );
  AOI22_X1 U3613 ( .A1(n6323), .A2(\dp/a_neg_mult_id_exe_int[2] ), .B1(n5184), 
        .B2(\dp/a_neg_mult_id_exe_int[3] ), .ZN(n3668) );
  AOI22_X1 U3614 ( .A1(n6322), .A2(\dp/a_mult_id_exe_int[3] ), .B1(
        \dp/mul_feedback_exe_mem_int[3] ), .B2(n5156), .ZN(n3669) );
  NAND2_X1 U3615 ( .A1(n3668), .A2(n3669), .ZN(n5840) );
  INV_X1 U3616 ( .A(n6704), .ZN(n3670) );
  AOI21_X1 U3617 ( .B1(n6703), .B2(n6303), .A(n6706), .ZN(n3671) );
  OAI21_X1 U3618 ( .B1(n6319), .B2(n3670), .A(n3671), .ZN(n6712) );
  AND2_X1 U3619 ( .A1(btb_cache_read_address[1]), .A2(
        btb_cache_read_address[0]), .ZN(\add_x_20/n28 ) );
  NOR2_X1 U3620 ( .A1(n5230), .A2(n365), .ZN(n3672) );
  AOI21_X1 U3621 ( .B1(\dp/ids/rp1[7] ), .B2(n4136), .A(n3672), .ZN(n6862) );
  NAND3_X1 U3622 ( .A1(n5088), .A2(n4266), .A3(cpu_is_reading), .ZN(n7188) );
  INV_X1 U3623 ( .A(n5351), .ZN(n3673) );
  NAND2_X1 U3624 ( .A1(n5352), .A2(n3673), .ZN(n3674) );
  OAI21_X1 U3625 ( .B1(n5622), .B2(n5344), .A(n3912), .ZN(n3675) );
  OAI221_X1 U3626 ( .B1(n5347), .B2(n4799), .C1(n5347), .C2(n3674), .A(n3675), 
        .ZN(\ctrl_u/n557 ) );
  AND2_X1 U3627 ( .A1(\ctrl_u/curr_exe[12] ), .A2(n5667), .ZN(n3676) );
  OAI221_X1 U3628 ( .B1(n3676), .B2(n7340), .C1(n3676), .C2(
        \ctrl_u/curr_mem_12 ), .A(rst_mem_wb_regs), .ZN(\ctrl_u/n468 ) );
  INV_X1 U3629 ( .A(n5534), .ZN(n3677) );
  INV_X1 U3630 ( .A(n5577), .ZN(n3678) );
  AOI21_X1 U3631 ( .B1(n7264), .B2(n3678), .A(n5578), .ZN(n3679) );
  NOR2_X1 U3632 ( .A1(instr_if[31]), .A2(n5567), .ZN(n3680) );
  OAI21_X1 U3633 ( .B1(n5550), .B2(n3680), .A(n5502), .ZN(n3681) );
  OAI211_X1 U3634 ( .C1(n5501), .C2(n3677), .A(n3679), .B(n3681), .ZN(n3682)
         );
  AOI22_X1 U3635 ( .A1(\ctrl_u/curr_id[40] ), .A2(n3941), .B1(n5641), .B2(
        n3682), .ZN(\ctrl_u/n245 ) );
  OAI21_X1 U3636 ( .B1(\ctrl_u/n73 ), .B2(n5599), .A(n5598), .ZN(\ctrl_u/n551 ) );
  AOI22_X1 U3637 ( .A1(\dp/a_neg_mult_id_exe_int[31] ), .A2(n5126), .B1(n6410), 
        .B2(n5194), .ZN(n1444) );
  INV_X1 U3638 ( .A(n5201), .ZN(n3683) );
  NAND2_X1 U3639 ( .A1(\dp/a_mult_id_exe_int[2] ), .A2(n3876), .ZN(n3684) );
  OAI21_X1 U3640 ( .B1(n3683), .B2(n6884), .A(n3684), .ZN(n2944) );
  NAND2_X1 U3641 ( .A1(n4141), .A2(n3956), .ZN(n3685) );
  NAND2_X1 U3642 ( .A1(n4393), .A2(n3896), .ZN(n3686) );
  OAI211_X1 U3643 ( .C1(n7042), .C2(n4820), .A(n3685), .B(n3686), .ZN(n2713)
         );
  NAND2_X1 U3644 ( .A1(\dp/ids/rp2[20] ), .A2(n3880), .ZN(n3687) );
  NAND2_X1 U3645 ( .A1(\dp/b_adder_id_exe_int[20] ), .A2(n5206), .ZN(n3688) );
  NAND4_X1 U3646 ( .A1(n6993), .A2(n6987), .A3(n3687), .A4(n3688), .ZN(n2665)
         );
  INV_X1 U3647 ( .A(n4863), .ZN(n3689) );
  NOR3_X1 U3648 ( .A1(n4902), .A2(n5029), .A3(n3689), .ZN(n4861) );
  INV_X1 U3649 ( .A(n5060), .ZN(n3690) );
  NAND3_X1 U3650 ( .A1(n4751), .A2(n3863), .A3(n3690), .ZN(n3691) );
  OAI211_X1 U3651 ( .C1(\intadd_1/n56 ), .C2(n4757), .A(\intadd_1/n57 ), .B(
        n3691), .ZN(n4753) );
  AOI22_X1 U3652 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/a_shiftn[42] ), .B1(
        n3946), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[43] ), .ZN(n3692) );
  NAND2_X1 U3653 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[43] ), .A2(n3945), .ZN(
        n3693) );
  OAI21_X1 U3654 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[43] ), .A(n3693), 
        .ZN(n3694) );
  AOI21_X1 U3655 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[42] ), 
        .A(n3694), .ZN(n3695) );
  NAND2_X1 U3656 ( .A1(n3692), .A2(n3695), .ZN(n6245) );
  AOI22_X1 U3657 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[45] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[45] ), .ZN(n3696) );
  AOI22_X1 U3658 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[44] ), .B1(
        \dp/mul_feedback_exe_mem_int[45] ), .B2(n5186), .ZN(n3697) );
  NAND2_X1 U3659 ( .A1(n3696), .A2(n3697), .ZN(n6248) );
  AOI22_X1 U3660 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[53] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[53] ), .ZN(n3698) );
  AOI22_X1 U3661 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[52] ), .B1(
        \dp/mul_feedback_exe_mem_int[53] ), .B2(n5186), .ZN(n3699) );
  NAND2_X1 U3662 ( .A1(n3698), .A2(n3699), .ZN(n6278) );
  AOI22_X1 U3663 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[55] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[55] ), .ZN(n3700) );
  AOI22_X1 U3664 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[54] ), .B1(
        \dp/mul_feedback_exe_mem_int[55] ), .B2(n5186), .ZN(n3701) );
  NAND2_X1 U3665 ( .A1(n3700), .A2(n3701), .ZN(n6285) );
  AOI22_X1 U3666 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[62] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[62] ), .ZN(n3702) );
  AOI22_X1 U3667 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[61] ), .B1(
        \dp/mul_feedback_exe_mem_int[62] ), .B2(n5186), .ZN(n3703) );
  NAND2_X1 U3668 ( .A1(n3702), .A2(n3703), .ZN(n6304) );
  INV_X1 U3669 ( .A(wp_data[2]), .ZN(n3704) );
  OAI22_X1 U3670 ( .A1(n5171), .A2(n3704), .B1(n5173), .B2(n4087), .ZN(n7247)
         );
  AND3_X1 U3671 ( .A1(n5239), .A2(\ctrl_u/curr_exe_40 ), .A3(
        \ctrl_u/curr_mem[3] ), .ZN(n4737) );
  AOI22_X1 U3672 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[28] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[29] ), .ZN(n3705) );
  AOI22_X1 U3673 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[29] ), .B1(
        \dp/mul_feedback_exe_mem_int[29] ), .B2(n5186), .ZN(n3706) );
  NAND2_X1 U3674 ( .A1(n3705), .A2(n3706), .ZN(n6118) );
  AOI222_X1 U3675 ( .A1(n5170), .A2(n4295), .B1(n4016), .B2(n4064), .C1(n5284), 
        .C2(n4043), .ZN(n3707) );
  INV_X1 U3676 ( .A(n3707), .ZN(n6096) );
  NAND2_X1 U3677 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[21] ), .A2(n6326), 
        .ZN(n3708) );
  NAND3_X1 U3678 ( .A1(n3708), .A2(n6025), .A3(n6026), .ZN(n6029) );
  AOI22_X1 U3679 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[15] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[16] ), .ZN(n3709) );
  AOI22_X1 U3680 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[16] ), .B1(
        \dp/mul_feedback_exe_mem_int[16] ), .B2(n5186), .ZN(n3710) );
  NAND2_X1 U3681 ( .A1(n3709), .A2(n3710), .ZN(n5756) );
  NAND2_X1 U3682 ( .A1(\dp/exs/alu_unit/mult/neg_ax2_shiftn[11] ), .A2(n6326), 
        .ZN(n3711) );
  AOI22_X1 U3683 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/ax2_shiftn[11] ), 
        .B1(n3945), .B2(\dp/exs/alu_unit/mult/ax2_shiftn[12] ), .ZN(n3712) );
  AOI21_X1 U3684 ( .B1(\dp/exs/alu_unit/mult/neg_ax2_shiftn[12] ), .B2(n3946), 
        .A(n5740), .ZN(n3713) );
  NAND3_X1 U3685 ( .A1(n3711), .A2(n3712), .A3(n3713), .ZN(n5922) );
  AOI22_X1 U3686 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[7] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[8] ), .ZN(n3714) );
  AOI22_X1 U3687 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[8] ), .B1(
        \dp/mul_feedback_exe_mem_int[8] ), .B2(n5156), .ZN(n3715) );
  NAND2_X1 U3688 ( .A1(n3714), .A2(n3715), .ZN(n5897) );
  INV_X1 U3689 ( .A(\intadd_1/n154 ), .ZN(n3716) );
  NOR2_X1 U3690 ( .A1(\intadd_1/n153 ), .A2(n3716), .ZN(n3717) );
  INV_X1 U3691 ( .A(\intadd_1/n159 ), .ZN(n3718) );
  AOI21_X1 U3692 ( .B1(\intadd_1/n160 ), .B2(\intadd_1/n196 ), .A(n3718), .ZN(
        n3719) );
  XNOR2_X1 U3693 ( .A(n3717), .B(n3719), .ZN(n4995) );
  AOI22_X1 U3694 ( .A1(n6298), .A2(\dp/exs/alu_unit/mult/a_shiftn[2] ), .B1(
        n5187), .B2(\dp/exs/alu_unit/mult/ax2_shiftn[4] ), .ZN(n3720) );
  AOI21_X1 U3695 ( .B1(\dp/exs/alu_unit/mult/neg_ax2_shiftn[4] ), .B2(n5188), 
        .A(n5702), .ZN(n3721) );
  NAND2_X1 U3696 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[2] ), .A2(n5154), 
        .ZN(n3722) );
  NAND3_X1 U3697 ( .A1(n3722), .A2(n3720), .A3(n3721), .ZN(n5841) );
  INV_X1 U3698 ( .A(n6514), .ZN(n3723) );
  INV_X1 U3699 ( .A(n6519), .ZN(n3724) );
  AOI21_X1 U3700 ( .B1(n6518), .B2(n6524), .A(n3724), .ZN(n3725) );
  NAND2_X1 U3701 ( .A1(n6219), .A2(n6512), .ZN(n3726) );
  OAI211_X1 U3702 ( .C1(n6315), .C2(n3723), .A(n3725), .B(n3726), .ZN(n6563)
         );
  OR2_X1 U3703 ( .A1(n6267), .A2(n6268), .ZN(n6598) );
  AOI21_X1 U3704 ( .B1(n5075), .B2(n5073), .A(n5041), .ZN(n3727) );
  XOR2_X1 U3705 ( .A(n4210), .B(\intadd_2/A[4] ), .Z(n3728) );
  XNOR2_X1 U3706 ( .A(n3727), .B(n3728), .ZN(\intadd_2/SUM[4] ) );
  AOI21_X1 U3707 ( .B1(n4032), .B2(n4829), .A(n4827), .ZN(n3729) );
  XOR2_X1 U3708 ( .A(\intadd_2/B[20] ), .B(n3866), .Z(n3730) );
  XNOR2_X1 U3709 ( .A(n3729), .B(n3730), .ZN(\intadd_2/SUM[20] ) );
  INV_X1 U3710 ( .A(n5349), .ZN(n3731) );
  OAI21_X1 U3711 ( .B1(n5164), .B2(n5350), .A(n3731), .ZN(n5355) );
  AOI21_X1 U3712 ( .B1(\intadd_2/n17 ), .B2(n4931), .A(n4929), .ZN(n3732) );
  XOR2_X1 U3713 ( .A(\intadd_2/B[14] ), .B(n4205), .Z(n3733) );
  XNOR2_X1 U3714 ( .A(n3732), .B(n3733), .ZN(\intadd_2/SUM[14] ) );
  INV_X1 U3715 ( .A(n4990), .ZN(n3734) );
  AOI21_X1 U3716 ( .B1(n4991), .B2(n5931), .A(n3734), .ZN(n3735) );
  XNOR2_X1 U3717 ( .A(n5940), .B(n5939), .ZN(n3736) );
  XNOR2_X1 U3718 ( .A(n3736), .B(n3735), .ZN(n3737) );
  NAND3_X1 U3719 ( .A1(n5012), .A2(\intadd_1/B[13] ), .A3(n3952), .ZN(n3738)
         );
  AOI21_X1 U3720 ( .B1(n5012), .B2(n7069), .A(\intadd_1/B[13] ), .ZN(n3739) );
  OAI21_X1 U3721 ( .B1(n3940), .B2(n5012), .A(n3739), .ZN(n3740) );
  OAI211_X1 U3722 ( .C1(\intadd_1/SUM[13] ), .C2(n7066), .A(n3738), .B(n3740), 
        .ZN(n3741) );
  AOI21_X1 U3723 ( .B1(\dp/exs/alu_unit/shifter_out[14] ), .B2(n3954), .A(
        n3741), .ZN(n3742) );
  OAI21_X1 U3724 ( .B1(n6027), .B2(n3737), .A(n3742), .ZN(n6437) );
  INV_X1 U3725 ( .A(n6701), .ZN(n3743) );
  AOI21_X1 U3726 ( .B1(n6693), .B2(n3743), .A(n6692), .ZN(n3744) );
  NAND2_X1 U3727 ( .A1(n6691), .A2(n6690), .ZN(n3745) );
  XOR2_X1 U3728 ( .A(n3744), .B(n3745), .Z(n6694) );
  NAND2_X1 U3729 ( .A1(n4136), .A2(\dp/ids/rp1[1] ), .ZN(n6889) );
  INV_X1 U3730 ( .A(\dp/ids/rp2[3] ), .ZN(n7050) );
  NAND2_X1 U3731 ( .A1(n5069), .A2(\intadd_1/n28 ), .ZN(n3746) );
  NAND3_X1 U3732 ( .A1(n3746), .A2(n5049), .A3(n5050), .ZN(n3747) );
  NAND2_X1 U3733 ( .A1(n5050), .A2(n4322), .ZN(n3748) );
  NAND3_X1 U3734 ( .A1(n3748), .A2(n5335), .A3(n3747), .ZN(n7092) );
  OAI22_X1 U3735 ( .A1(btb_cache_read_address[0]), .A2(n7105), .B1(n7109), 
        .B2(btb_cache_rw_address[0]), .ZN(n3749) );
  INV_X1 U3736 ( .A(n3749), .ZN(n4002) );
  AOI22_X1 U3737 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[18] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[18] ), .ZN(n3750) );
  INV_X1 U3738 ( .A(n3750), .ZN(wp_data[18]) );
  AOI22_X1 U3739 ( .A1(n4336), .A2(n4090), .B1(n5228), .B2(n4282), .ZN(
        wp_data[25]) );
  INV_X1 U3740 ( .A(n7340), .ZN(n3751) );
  AOI221_X1 U3741 ( .B1(\ctrl_u/curr_mem[2] ), .B2(n3751), .C1(wp_en), .C2(
        n7340), .A(n5229), .ZN(\ctrl_u/n483 ) );
  AND2_X1 U3742 ( .A1(\ctrl_u/curr_exe[13] ), .A2(n5667), .ZN(n3752) );
  OAI221_X1 U3743 ( .B1(n3752), .B2(n7340), .C1(n3752), .C2(wr_mem), .A(
        rst_mem_wb_regs), .ZN(\ctrl_u/n467 ) );
  INV_X1 U3744 ( .A(n5511), .ZN(n3753) );
  NAND3_X1 U3745 ( .A1(n5540), .A2(n5518), .A3(n5530), .ZN(n3754) );
  NAND3_X1 U3746 ( .A1(n5624), .A2(n5513), .A3(n3754), .ZN(n3755) );
  AOI211_X1 U3747 ( .C1(instr_if[27]), .C2(n3753), .A(n5575), .B(n3755), .ZN(
        n3756) );
  OAI22_X1 U3748 ( .A1(n5182), .A2(n4601), .B1(n3756), .B2(n5653), .ZN(
        \ctrl_u/n524 ) );
  OAI21_X1 U3749 ( .B1(\ctrl_u/n74 ), .B2(n5599), .A(n5598), .ZN(\ctrl_u/n552 ) );
  INV_X1 U3750 ( .A(n5618), .ZN(n3757) );
  OAI211_X1 U3751 ( .C1(n5617), .C2(n3757), .A(n5655), .B(n4237), .ZN(n3758)
         );
  NAND2_X1 U3752 ( .A1(n5670), .A2(n3758), .ZN(n3759) );
  NOR2_X1 U3753 ( .A1(n3757), .A2(n3759), .ZN(n3760) );
  AOI211_X1 U3754 ( .C1(\ctrl_u/n83 ), .C2(n3759), .A(n5619), .B(n3760), .ZN(
        \ctrl_u/n69 ) );
  AOI211_X1 U3755 ( .C1(n3936), .C2(\dp/pc_plus4_out_if_int[22] ), .A(n5018), 
        .B(n4133), .ZN(n3761) );
  AOI22_X1 U3756 ( .A1(btb_cache_read_address[22]), .A2(n5193), .B1(
        \dp/ifs/pc_btb[22] ), .B2(n3931), .ZN(n3762) );
  NAND2_X1 U3757 ( .A1(n4893), .A2(n3883), .ZN(n3763) );
  NAND3_X1 U3758 ( .A1(n3763), .A2(n3761), .A3(n3762), .ZN(n2535) );
  AOI22_X1 U3759 ( .A1(\dp/a_neg_mult_id_exe_int[10] ), .A2(n5127), .B1(n4888), 
        .B2(n7097), .ZN(n1466) );
  AOI22_X1 U3760 ( .A1(\dp/ids/rp2[31] ), .A2(n5214), .B1(
        \dp/id_exe_regs/b_mult_reg/q[30] ), .B2(n3897), .ZN(n3764) );
  NAND2_X1 U3761 ( .A1(n6963), .A2(n3764), .ZN(n2686) );
  NAND2_X1 U3762 ( .A1(\dp/ids/rp2[19] ), .A2(n3881), .ZN(n3765) );
  NAND2_X1 U3763 ( .A1(\dp/b_adder_id_exe_int[19] ), .A2(n5207), .ZN(n3766) );
  NAND4_X1 U3764 ( .A1(n6993), .A2(n6989), .A3(n3765), .A4(n3766), .ZN(n2666)
         );
  INV_X1 U3765 ( .A(n5200), .ZN(n3767) );
  NAND2_X1 U3766 ( .A1(\dp/b10_1_mult_id_exe_int[1] ), .A2(n3878), .ZN(n3768)
         );
  OAI21_X1 U3767 ( .B1(n3767), .B2(n7061), .A(n3768), .ZN(n2723) );
  AOI22_X1 U3768 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[30] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[30] ), .ZN(n3769) );
  AOI22_X1 U3769 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[29] ), .B1(
        \dp/mul_feedback_exe_mem_int[30] ), .B2(n5186), .ZN(n3770) );
  NAND2_X1 U3770 ( .A1(n3769), .A2(n3770), .ZN(n6140) );
  AOI22_X1 U3771 ( .A1(n5189), .A2(\dp/exs/alu_unit/mult/a_shiftn[35] ), .B1(
        n3945), .B2(\dp/exs/alu_unit/mult/a_shiftn[36] ), .ZN(n3771) );
  NAND2_X1 U3772 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[36] ), .A2(n3946), 
        .ZN(n3772) );
  OAI21_X1 U3773 ( .B1(n5169), .B2(\dp/a_mult_id_exe_int[36] ), .A(n3772), 
        .ZN(n3773) );
  AOI21_X1 U3774 ( .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[35] ), 
        .A(n3773), .ZN(n3774) );
  NAND2_X1 U3775 ( .A1(n3771), .A2(n3774), .ZN(n6211) );
  INV_X1 U3776 ( .A(n5073), .ZN(n3775) );
  AOI22_X1 U3777 ( .A1(\dp/npc_id_exe_int[7] ), .A2(n4130), .B1(n5072), .B2(
        n3775), .ZN(n5040) );
  NOR2_X1 U3778 ( .A1(n5494), .A2(instr_if[30]), .ZN(n3776) );
  AOI211_X1 U3779 ( .C1(n5494), .C2(instr_if[30]), .A(n5649), .B(n3776), .ZN(
        n5604) );
  AOI21_X1 U3780 ( .B1(\intadd_1/n68 ), .B2(\intadd_1/n89 ), .A(\intadd_1/n69 ), .ZN(n3777) );
  NAND2_X1 U3781 ( .A1(\intadd_1/n65 ), .A2(n5059), .ZN(n3778) );
  XOR2_X1 U3782 ( .A(n3777), .B(n3778), .Z(\intadd_1/SUM[19] ) );
  NOR2_X1 U3783 ( .A1(n4746), .A2(n4131), .ZN(n3779) );
  AOI21_X1 U3784 ( .B1(n4211), .B2(n4137), .A(n3779), .ZN(n4745) );
  AOI22_X1 U3785 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[27] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[28] ), .ZN(n3780) );
  AOI22_X1 U3786 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[28] ), .B1(
        \dp/mul_feedback_exe_mem_int[28] ), .B2(n5186), .ZN(n3781) );
  NAND2_X1 U3787 ( .A1(n3780), .A2(n3781), .ZN(n6135) );
  NAND2_X1 U3788 ( .A1(n5170), .A2(n4307), .ZN(n3782) );
  INV_X1 U3789 ( .A(n4041), .ZN(n3783) );
  OAI21_X1 U3790 ( .B1(n4024), .B2(n4062), .A(n3783), .ZN(n3784) );
  OAI211_X1 U3791 ( .C1(n5273), .C2(wp_data[25]), .A(n3782), .B(n3784), .ZN(
        n6065) );
  INV_X1 U3792 ( .A(n5077), .ZN(n3785) );
  NOR2_X1 U3793 ( .A1(n5068), .A2(n3785), .ZN(n4206) );
  AOI22_X1 U3794 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[14] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[15] ), .ZN(n3786) );
  AOI22_X1 U3795 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[15] ), .B1(
        \dp/mul_feedback_exe_mem_int[15] ), .B2(n5186), .ZN(n3787) );
  NAND2_X1 U3796 ( .A1(n3786), .A2(n3787), .ZN(n5942) );
  AOI22_X1 U3797 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[12] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[13] ), .ZN(n3788) );
  AOI22_X1 U3798 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[13] ), .B1(
        \dp/mul_feedback_exe_mem_int[13] ), .B2(n5186), .ZN(n3789) );
  NAND2_X1 U3799 ( .A1(n3788), .A2(n3789), .ZN(n5929) );
  AOI22_X1 U3800 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[10] ), .B1(n3939), 
        .B2(\dp/a_neg_mult_id_exe_int[11] ), .ZN(n3790) );
  AOI22_X1 U3801 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[11] ), .B1(
        \dp/mul_feedback_exe_mem_int[11] ), .B2(n5186), .ZN(n3791) );
  NAND2_X1 U3802 ( .A1(n3790), .A2(n3791), .ZN(n5921) );
  AOI22_X1 U3803 ( .A1(n5156), .A2(\dp/mul_feedback_exe_mem_int[7] ), .B1(
        \dp/a_neg_mult_id_exe_int[6] ), .B2(n3919), .ZN(n3792) );
  NAND3_X1 U3804 ( .A1(n5727), .A2(n5728), .A3(n3792), .ZN(n5885) );
  INV_X1 U3805 ( .A(\intadd_1/n149 ), .ZN(n3793) );
  NOR2_X1 U3806 ( .A1(\intadd_1/n148 ), .A2(n3793), .ZN(n3794) );
  XNOR2_X1 U3807 ( .A(\intadd_1/n150 ), .B(n3794), .ZN(\intadd_1/SUM[5] ) );
  OR2_X1 U3808 ( .A1(n6196), .A2(n6197), .ZN(n6478) );
  OR2_X1 U3809 ( .A1(n6217), .A2(n6218), .ZN(n6519) );
  OR2_X1 U3810 ( .A1(n6238), .A2(n6239), .ZN(n6533) );
  AOI21_X1 U3811 ( .B1(n6614), .B2(n6615), .A(n6613), .ZN(n3795) );
  INV_X1 U3812 ( .A(n3795), .ZN(n4919) );
  INV_X1 U3813 ( .A(n6643), .ZN(n3796) );
  INV_X1 U3814 ( .A(n6287), .ZN(n3797) );
  NOR2_X1 U3815 ( .A1(n6662), .A2(n3797), .ZN(n3798) );
  AOI211_X1 U3816 ( .C1(n6676), .C2(n6673), .A(n3798), .B(n6677), .ZN(n3799)
         );
  NAND2_X1 U3817 ( .A1(n6317), .A2(n6625), .ZN(n3800) );
  OAI211_X1 U3818 ( .C1(n6282), .C2(n3796), .A(n3799), .B(n3800), .ZN(n6682)
         );
  INV_X1 U3819 ( .A(\dp/exs/alu_unit/mult/a_shiftn[62] ), .ZN(n3801) );
  AOI22_X1 U3820 ( .A1(n5188), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[63] ), 
        .B1(n6326), .B2(\dp/exs/alu_unit/mult/neg_a_shiftn[62] ), .ZN(n3802)
         );
  AOI22_X1 U3821 ( .A1(n3945), .A2(\dp/exs/alu_unit/mult/a_shiftn[63] ), .B1(
        n6327), .B2(n4493), .ZN(n3803) );
  OAI211_X1 U3822 ( .C1(n6328), .C2(n3801), .A(n3802), .B(n3803), .ZN(n6329)
         );
  AOI21_X1 U3823 ( .B1(n4795), .B2(n4802), .A(n4320), .ZN(n3804) );
  NAND3_X1 U3824 ( .A1(n4732), .A2(n4731), .A3(n4775), .ZN(n3805) );
  OAI21_X1 U3825 ( .B1(n4256), .B2(n3804), .A(n3805), .ZN(n3806) );
  INV_X1 U3826 ( .A(n3806), .ZN(\intadd_1/n28 ) );
  NAND3_X1 U3827 ( .A1(ram_update), .A2(n4371), .A3(wr_mem), .ZN(n3807) );
  NOR2_X1 U3828 ( .A1(\mc/currstate[1] ), .A2(n3807), .ZN(n5809) );
  NAND2_X1 U3829 ( .A1(n4136), .A2(\dp/ids/rp1[0] ), .ZN(n6894) );
  INV_X1 U3830 ( .A(\dp/ids/rp2[2] ), .ZN(n7103) );
  AOI21_X1 U3831 ( .B1(n7298), .B2(\ctrl_u/curr_exe[17] ), .A(n7442), .ZN(
        n7426) );
  AOI22_X1 U3832 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[0] ), .B1(n5228), 
        .B2(\dp/cache_data_mem_wb_int[0] ), .ZN(n3808) );
  INV_X1 U3833 ( .A(n3808), .ZN(wp_data[0]) );
  AOI22_X1 U3834 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[1] ), .B1(n5228), 
        .B2(\dp/cache_data_mem_wb_int[1] ), .ZN(n3809) );
  INV_X1 U3835 ( .A(n3809), .ZN(wp_data[1]) );
  AOI22_X1 U3836 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[2] ), .B1(n5228), 
        .B2(\dp/cache_data_mem_wb_int[2] ), .ZN(n3810) );
  INV_X1 U3837 ( .A(n3810), .ZN(wp_data[2]) );
  AOI22_X1 U3838 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[3] ), .B1(n5228), 
        .B2(\dp/cache_data_mem_wb_int[3] ), .ZN(n3811) );
  INV_X1 U3839 ( .A(n3811), .ZN(wp_data[3]) );
  AOI22_X1 U3840 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[4] ), .B1(n5228), 
        .B2(\dp/cache_data_mem_wb_int[4] ), .ZN(n3812) );
  INV_X1 U3841 ( .A(n3812), .ZN(wp_data[4]) );
  AOI22_X1 U3842 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[5] ), .B1(n5228), 
        .B2(\dp/cache_data_mem_wb_int[5] ), .ZN(n3813) );
  INV_X1 U3843 ( .A(n3813), .ZN(wp_data[5]) );
  AOI22_X1 U3844 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[6] ), .B1(n5228), 
        .B2(\dp/cache_data_mem_wb_int[6] ), .ZN(n3814) );
  INV_X1 U3845 ( .A(n3814), .ZN(wp_data[6]) );
  AOI22_X1 U3846 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[7] ), .B1(n5228), 
        .B2(\dp/cache_data_mem_wb_int[7] ), .ZN(n3815) );
  INV_X1 U3847 ( .A(n3815), .ZN(wp_data[7]) );
  AOI22_X1 U3848 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[8] ), .B1(n5228), 
        .B2(\dp/cache_data_mem_wb_int[8] ), .ZN(n3816) );
  INV_X1 U3849 ( .A(n3816), .ZN(wp_data[8]) );
  AOI22_X1 U3850 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[9] ), .B1(n5228), 
        .B2(\dp/cache_data_mem_wb_int[9] ), .ZN(n3817) );
  INV_X1 U3851 ( .A(n3817), .ZN(wp_data[9]) );
  AOI22_X1 U3852 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[10] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[10] ), .ZN(n3818) );
  INV_X1 U3853 ( .A(n3818), .ZN(wp_data[10]) );
  AOI22_X1 U3854 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[11] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[11] ), .ZN(n3819) );
  INV_X1 U3855 ( .A(n3819), .ZN(wp_data[11]) );
  AOI22_X1 U3856 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[12] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[12] ), .ZN(n3820) );
  INV_X1 U3857 ( .A(n3820), .ZN(wp_data[12]) );
  AOI22_X1 U3858 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[13] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[13] ), .ZN(n3821) );
  INV_X1 U3859 ( .A(n3821), .ZN(wp_data[13]) );
  AOI22_X1 U3860 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[14] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[14] ), .ZN(n3822) );
  INV_X1 U3861 ( .A(n3822), .ZN(wp_data[14]) );
  AOI22_X1 U3862 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[15] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[15] ), .ZN(n3823) );
  INV_X1 U3863 ( .A(n3823), .ZN(wp_data[15]) );
  AOI22_X1 U3864 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[16] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[16] ), .ZN(n3824) );
  INV_X1 U3865 ( .A(n3824), .ZN(wp_data[16]) );
  AOI22_X1 U3866 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[17] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[17] ), .ZN(n3825) );
  INV_X1 U3867 ( .A(n3825), .ZN(wp_data[17]) );
  AOI22_X1 U3868 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[19] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[19] ), .ZN(n3826) );
  INV_X1 U3869 ( .A(n3826), .ZN(wp_data[19]) );
  AOI22_X1 U3870 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[20] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[20] ), .ZN(n3827) );
  INV_X1 U3871 ( .A(n3827), .ZN(wp_data[20]) );
  AOI22_X1 U3872 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[21] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[21] ), .ZN(n3828) );
  INV_X1 U3873 ( .A(n3828), .ZN(wp_data[21]) );
  AOI22_X1 U3874 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[22] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[22] ), .ZN(n3829) );
  INV_X1 U3875 ( .A(n3829), .ZN(wp_data[22]) );
  AOI22_X1 U3876 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[23] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[23] ), .ZN(n3830) );
  INV_X1 U3877 ( .A(n3830), .ZN(wp_data[23]) );
  AOI22_X1 U3878 ( .A1(n4336), .A2(n4112), .B1(n5228), .B2(n4283), .ZN(
        wp_data[24]) );
  AOI22_X1 U3879 ( .A1(n4336), .A2(n4091), .B1(n5228), .B2(n4281), .ZN(
        wp_data[26]) );
  AOI22_X1 U3880 ( .A1(n4336), .A2(n4092), .B1(n5228), .B2(n4280), .ZN(
        wp_data[27]) );
  AOI22_X1 U3881 ( .A1(n4336), .A2(n4093), .B1(n5228), .B2(n4279), .ZN(
        wp_data[28]) );
  AOI22_X1 U3882 ( .A1(n4336), .A2(n4094), .B1(n5228), .B2(n4278), .ZN(
        wp_data[29]) );
  AOI22_X1 U3883 ( .A1(n4336), .A2(n7496), .B1(n5228), .B2(n4277), .ZN(
        wp_data[30]) );
  AOI22_X1 U3884 ( .A1(n4336), .A2(\dp/alu_out_low_mem_wb_int[31] ), .B1(n5228), .B2(\dp/cache_data_mem_wb_int[31] ), .ZN(n3831) );
  INV_X1 U3885 ( .A(n3831), .ZN(wp_data[31]) );
  NOR3_X1 U3886 ( .A1(n3981), .A2(n7340), .A3(n5824), .ZN(
        btb_cache_update_line) );
  INV_X1 U3887 ( .A(n7340), .ZN(n3832) );
  OAI221_X1 U3888 ( .B1(n7340), .B2(\ctrl_u/curr_mem[1] ), .C1(n3832), .C2(
        n5228), .A(rst_mem_wb_regs), .ZN(\ctrl_u/n484 ) );
  AOI21_X1 U3889 ( .B1(n5568), .B2(n5572), .A(n5584), .ZN(n3833) );
  AOI21_X1 U3890 ( .B1(\ctrl_u/curr_id[39] ), .B2(n3941), .A(n3833), .ZN(n3834) );
  NAND2_X1 U3891 ( .A1(n5547), .A2(n3834), .ZN(\ctrl_u/n523 ) );
  INV_X1 U3892 ( .A(n7340), .ZN(n3835) );
  OAI221_X1 U3893 ( .B1(n7340), .B2(\ctrl_u/curr_mem[0] ), .C1(n3835), .C2(
        hilo_wr_en), .A(rst_mem_wb_regs), .ZN(\ctrl_u/n486 ) );
  OR2_X1 U3894 ( .A1(\ctrl_u/curr_wb[3] ), .A2(n5670), .ZN(n3836) );
  AOI221_X1 U3895 ( .B1(n7340), .B2(n3836), .C1(\ctrl_u/curr_mem[3] ), .C2(
        n3836), .A(n5229), .ZN(\ctrl_u/n481 ) );
  AND2_X1 U3896 ( .A1(\ctrl_u/curr_exe[14] ), .A2(n5667), .ZN(n3837) );
  OAI221_X1 U3897 ( .B1(n3837), .B2(cpu_is_reading), .C1(n3837), .C2(n7340), 
        .A(rst_mem_wb_regs), .ZN(\ctrl_u/n465 ) );
  NOR2_X1 U3898 ( .A1(n5162), .A2(n5350), .ZN(n3838) );
  NOR2_X1 U3899 ( .A1(n5355), .A2(n3838), .ZN(n3839) );
  INV_X1 U3900 ( .A(n5149), .ZN(n3840) );
  NAND2_X1 U3901 ( .A1(n5354), .A2(n3840), .ZN(n3841) );
  OAI22_X1 U3902 ( .A1(n5348), .A2(n3841), .B1(n3839), .B2(n3840), .ZN(
        \ctrl_u/n504 ) );
  NAND2_X1 U3903 ( .A1(n5624), .A2(n5625), .ZN(n3842) );
  INV_X1 U3904 ( .A(n5626), .ZN(n3843) );
  OAI221_X1 U3905 ( .B1(n5626), .B2(n3842), .C1(n3843), .C2(n4492), .A(n4815), 
        .ZN(\ctrl_u/n535 ) );
  OAI22_X1 U3906 ( .A1(n6694), .A2(n7062), .B1(n4204), .B2(n3938), .ZN(n2791)
         );
  AOI22_X1 U3907 ( .A1(\dp/ids/rp2[30] ), .A2(n5214), .B1(
        \dp/id_exe_regs/b_mult_reg/q[29] ), .B2(n3898), .ZN(n3844) );
  NAND2_X1 U3908 ( .A1(n6963), .A2(n3844), .ZN(n2687) );
  INV_X1 U3909 ( .A(n5215), .ZN(n3845) );
  AOI222_X1 U3910 ( .A1(n3845), .A2(\dp/ids/rp2[25] ), .B1(
        \dp/op_b_id_ex_int[25] ), .B2(n7100), .C1(n4409), .C2(n4107), .ZN(
        n3846) );
  INV_X1 U3911 ( .A(n3846), .ZN(n2731) );
  NAND2_X1 U3912 ( .A1(\dp/ids/rp2[18] ), .A2(n3881), .ZN(n3847) );
  NAND2_X1 U3913 ( .A1(\dp/b_adder_id_exe_int[18] ), .A2(n5208), .ZN(n3848) );
  NAND4_X1 U3914 ( .A1(n6993), .A2(n6992), .A3(n3847), .A4(n3848), .ZN(n2667)
         );
  INV_X1 U3915 ( .A(n5200), .ZN(n3849) );
  NAND2_X1 U3916 ( .A1(n4231), .A2(n3878), .ZN(n3850) );
  OAI21_X1 U3917 ( .B1(n3849), .B2(n7054), .A(n3850), .ZN(n2722) );
  INV_X1 U3918 ( .A(n7084), .ZN(n3851) );
  AOI22_X1 U3919 ( .A1(\dp/a_neg_mult_id_exe_int[0] ), .A2(n5126), .B1(n7097), 
        .B2(n3851), .ZN(n1493) );
  AOI22_X1 U3920 ( .A1(btb_cache_read_address[0]), .A2(n5193), .B1(
        \dp/ifs/pc_btb[0] ), .B2(n3895), .ZN(n3852) );
  AOI22_X1 U3921 ( .A1(n4892), .A2(n3884), .B1(n7107), .B2(n3926), .ZN(n3853)
         );
  NAND3_X1 U3922 ( .A1(n4002), .A2(n3852), .A3(n3853), .ZN(n2557) );
  XOR2_X1 U3923 ( .A(btb_cache_read_address[0]), .B(btb_cache_read_address[1]), 
        .Z(\dp/pc_plus4_out_if_int[1] ) );
  BUF_X1 U3924 ( .A(n4039), .Z(n3854) );
  BUF_X1 U3925 ( .A(n4923), .Z(n3855) );
  NOR2_X2 U3926 ( .A1(n7177), .A2(n3856), .ZN(n5581) );
  AND2_X1 U3927 ( .A1(n4816), .A2(\ctrl_u/if_stall ), .ZN(n3856) );
  AND2_X1 U3928 ( .A1(n4875), .A2(n5044), .ZN(n4054) );
  OR2_X1 U3929 ( .A1(n3927), .A2(n4856), .ZN(n3857) );
  BUF_X1 U3930 ( .A(n4968), .Z(n3858) );
  BUF_X1 U3931 ( .A(n3948), .Z(n3859) );
  INV_X1 U3932 ( .A(\intadd_1/n182 ), .ZN(n3860) );
  BUF_X1 U3933 ( .A(\intadd_1/n74 ), .Z(n3861) );
  BUF_X1 U3934 ( .A(\intadd_1/SUM[17] ), .Z(n3862) );
  INV_X1 U3935 ( .A(n4758), .ZN(n3863) );
  BUF_X1 U3936 ( .A(\intadd_1/SUM[28] ), .Z(n3864) );
  NOR2_X1 U3937 ( .A1(\intadd_1/n64 ), .A2(\intadd_1/n61 ), .ZN(\intadd_1/n59 ) );
  BUF_X2 U3938 ( .A(n7272), .Z(n3906) );
  NAND2_X1 U3939 ( .A1(n3932), .A2(n6721), .ZN(n3865) );
  BUF_X1 U3940 ( .A(n5176), .Z(n4052) );
  INV_X2 U3941 ( .A(n4052), .ZN(n4850) );
  BUF_X2 U3942 ( .A(n6323), .Z(n3943) );
  NAND2_X2 U3943 ( .A1(n7171), .A2(n6473), .ZN(n7058) );
  INV_X2 U3944 ( .A(n4228), .ZN(n5226) );
  BUF_X2 U3945 ( .A(n7100), .Z(n5129) );
  BUF_X2 U3946 ( .A(n7100), .Z(n5128) );
  AND2_X2 U3947 ( .A1(n3901), .A2(n4921), .ZN(n7097) );
  BUF_X4 U3948 ( .A(n7097), .Z(n5194) );
  OR2_X1 U3949 ( .A1(n5683), .A2(n593), .ZN(n5151) );
  NOR2_X2 U3950 ( .A1(n5683), .A2(n593), .ZN(n5184) );
  BUF_X4 U3951 ( .A(n5184), .Z(n3939) );
  BUF_X1 U3952 ( .A(n5168), .Z(n3900) );
  BUF_X4 U3953 ( .A(n3900), .Z(n5169) );
  INV_X2 U3954 ( .A(n3888), .ZN(n3893) );
  INV_X2 U3955 ( .A(n5138), .ZN(n4040) );
  BUF_X4 U3956 ( .A(n6719), .Z(n5196) );
  CLKBUF_X3 U3957 ( .A(n6756), .Z(n4057) );
  NAND2_X1 U3958 ( .A1(n7056), .A2(n6722), .ZN(n6756) );
  CLKBUF_X3 U3959 ( .A(n6756), .Z(n4056) );
  BUF_X2 U3960 ( .A(n5653), .Z(n3927) );
  BUF_X1 U3961 ( .A(n3944), .Z(n3930) );
  XOR2_X1 U3962 ( .A(n4257), .B(n4113), .Z(n3867) );
  NAND2_X1 U3963 ( .A1(n5044), .A2(btb_cache_update_line), .ZN(n3870) );
  NOR2_X2 U3964 ( .A1(\intadd_1/A[8] ), .A2(\intadd_1/B[8] ), .ZN(
        \intadd_1/n134 ) );
  OR2_X4 U3965 ( .A1(n5142), .A2(\ctrl_u/curr_exe_39 ), .ZN(n3922) );
  INV_X1 U3966 ( .A(n6701), .ZN(n3871) );
  NOR2_X2 U3967 ( .A1(n5140), .A2(n5141), .ZN(n5122) );
  BUF_X2 U3968 ( .A(n7272), .Z(n5140) );
  NAND2_X2 U3969 ( .A1(n4132), .A2(n4586), .ZN(n5618) );
  AND2_X1 U3970 ( .A1(n6311), .A2(n6310), .ZN(n3872) );
  AND4_X2 U3971 ( .A1(n4767), .A2(n4769), .A3(n4765), .A4(n4764), .ZN(n4989)
         );
  NAND2_X1 U3972 ( .A1(n5338), .A2(rst_mem_wb_regs), .ZN(n4968) );
  OR2_X2 U3973 ( .A1(n3981), .A2(n5824), .ZN(n5338) );
  OAI21_X2 U3974 ( .B1(n6177), .B2(\ctrl_u/curr_exe[20] ), .A(n6176), .ZN(
        n6182) );
  BUF_X4 U3975 ( .A(n7109), .Z(n3873) );
  BUF_X1 U3976 ( .A(n7060), .Z(n3874) );
  BUF_X1 U3977 ( .A(n7060), .Z(n3875) );
  INV_X2 U3978 ( .A(n5181), .ZN(n3935) );
  CLKBUF_X3 U3979 ( .A(n7272), .Z(n4024) );
  NOR2_X2 U3980 ( .A1(n5768), .A2(n4738), .ZN(n7272) );
  BUF_X1 U3981 ( .A(n7272), .Z(n5139) );
  AND3_X1 U3982 ( .A1(n4798), .A2(n4726), .A3(n5096), .ZN(n7253) );
  AND2_X1 U3983 ( .A1(n4726), .A2(n5096), .ZN(n5137) );
  INV_X2 U3984 ( .A(n3865), .ZN(n3876) );
  INV_X2 U3985 ( .A(n3865), .ZN(n3877) );
  INV_X2 U3986 ( .A(n3865), .ZN(n3878) );
  NAND2_X1 U3987 ( .A1(n6179), .A2(taken), .ZN(n7104) );
  OR2_X1 U3988 ( .A1(n4876), .A2(n4821), .ZN(n3882) );
  OR2_X2 U3989 ( .A1(n4876), .A2(n4821), .ZN(n5414) );
  AND2_X1 U3990 ( .A1(n6180), .A2(n6182), .ZN(n3883) );
  AND2_X2 U3991 ( .A1(n6180), .A2(n6182), .ZN(n3884) );
  INV_X1 U3992 ( .A(n3883), .ZN(n3885) );
  NAND2_X2 U3993 ( .A1(n6931), .A2(n6930), .ZN(n5215) );
  AND2_X1 U3994 ( .A1(n6311), .A2(n6310), .ZN(n3886) );
  INV_X1 U3995 ( .A(n7138), .ZN(n3887) );
  INV_X1 U3996 ( .A(n7138), .ZN(n3888) );
  INV_X1 U3997 ( .A(n3887), .ZN(n3889) );
  INV_X1 U3998 ( .A(n3887), .ZN(n3890) );
  INV_X1 U3999 ( .A(n3887), .ZN(n3891) );
  INV_X1 U4000 ( .A(n3887), .ZN(n3892) );
  OR2_X1 U4001 ( .A1(n7141), .A2(en_npc_id), .ZN(n7138) );
  AND2_X1 U4002 ( .A1(n4875), .A2(n5044), .ZN(n3894) );
  AND2_X1 U4003 ( .A1(n4875), .A2(n5044), .ZN(n3895) );
  NAND2_X1 U4004 ( .A1(n4664), .A2(n5023), .ZN(n3901) );
  NAND2_X1 U4005 ( .A1(n4664), .A2(n5023), .ZN(n3902) );
  NAND2_X2 U4006 ( .A1(n4664), .A2(n5023), .ZN(n7171) );
  NOR2_X1 U4007 ( .A1(n5139), .A2(n5141), .ZN(n3903) );
  NOR2_X2 U4008 ( .A1(n3906), .A2(n5141), .ZN(n5120) );
  NOR2_X2 U4009 ( .A1(n5139), .A2(n5141), .ZN(n5119) );
  INV_X1 U4010 ( .A(n4517), .ZN(n3904) );
  BUF_X4 U4011 ( .A(n7253), .Z(n3949) );
  AND2_X2 U4012 ( .A1(n5249), .A2(n5248), .ZN(n5116) );
  NOR2_X1 U4013 ( .A1(\intadd_1/A[18] ), .A2(\intadd_1/B[18] ), .ZN(
        \intadd_1/n74 ) );
  INV_X1 U4014 ( .A(\intadd_1/n198 ), .ZN(n3905) );
  NOR2_X1 U4015 ( .A1(\intadd_1/B[1] ), .A2(\intadd_1/A[1] ), .ZN(
        \intadd_1/n167 ) );
  AND4_X2 U4016 ( .A1(n4736), .A2(n4737), .A3(n3909), .A4(n4735), .ZN(n4232)
         );
  BUF_X1 U4017 ( .A(n7272), .Z(n5138) );
  XOR2_X1 U4018 ( .A(n4489), .B(rd_exemem[1]), .Z(n5265) );
  AND2_X2 U4019 ( .A1(n5098), .A2(n5097), .ZN(n5096) );
  CLKBUF_X1 U4020 ( .A(n7273), .Z(n3933) );
  NOR2_X1 U4021 ( .A1(\intadd_1/A[6] ), .A2(\intadd_1/B[6] ), .ZN(
        \intadd_1/n145 ) );
  BUF_X2 U4022 ( .A(n5325), .Z(n5118) );
  NOR2_X2 U4023 ( .A1(dcache_hit), .A2(wr_mem), .ZN(n5088) );
  NAND2_X1 U4024 ( .A1(n6098), .A2(n6099), .ZN(n3907) );
  BUF_X1 U4025 ( .A(n5919), .Z(n3908) );
  NAND3_X2 U4026 ( .A1(n4797), .A2(n4726), .A3(n5096), .ZN(n5123) );
  AOI21_X2 U4027 ( .B1(n5065), .B2(n5077), .A(n5066), .ZN(n5064) );
  BUF_X1 U4028 ( .A(n4960), .Z(n3909) );
  OR2_X2 U4029 ( .A1(\mc/currstate[1] ), .A2(n4371), .ZN(n3910) );
  NAND2_X4 U4030 ( .A1(n5137), .A2(n4797), .ZN(n5173) );
  INV_X1 U4031 ( .A(n4025), .ZN(n3912) );
  INV_X1 U4032 ( .A(n3906), .ZN(n3913) );
  OR2_X1 U4033 ( .A1(\intadd_1/A[12] ), .A2(\intadd_1/B[12] ), .ZN(n3914) );
  NAND2_X1 U4034 ( .A1(n4874), .A2(n4873), .ZN(n3915) );
  BUF_X1 U4035 ( .A(\intadd_1/n97 ), .Z(n3916) );
  BUF_X2 U4036 ( .A(n5135), .Z(n5170) );
  BUF_X1 U4037 ( .A(n6088), .Z(n3917) );
  BUF_X1 U4038 ( .A(n5911), .Z(n3918) );
  BUF_X4 U4039 ( .A(n3943), .Z(n3919) );
  NOR2_X2 U4040 ( .A1(n5712), .A2(n5681), .ZN(n6323) );
  BUF_X1 U4041 ( .A(n5143), .Z(n3920) );
  BUF_X4 U4042 ( .A(n5187), .Z(n3945) );
  XNOR2_X1 U4043 ( .A(n3921), .B(n6481), .ZN(n6482) );
  AND2_X1 U4044 ( .A1(n6478), .A2(n6477), .ZN(n3921) );
  BUF_X1 U4045 ( .A(n5005), .Z(n3923) );
  AND4_X1 U4046 ( .A1(n4799), .A2(n5234), .A3(n4238), .A4(n5618), .ZN(n3924)
         );
  INV_X4 U4047 ( .A(n7177), .ZN(n5177) );
  CLKBUF_X3 U4048 ( .A(n5581), .Z(n5182) );
  BUF_X2 U4049 ( .A(n7186), .Z(n5179) );
  AND2_X2 U4050 ( .A1(n3932), .A2(n4914), .ZN(n7056) );
  INV_X4 U4051 ( .A(n3951), .ZN(n5185) );
  AND2_X2 U4052 ( .A1(n5150), .A2(n3899), .ZN(n5156) );
  BUF_X2 U4053 ( .A(n4816), .Z(n3929) );
  AND4_X2 U4054 ( .A1(n5234), .A2(n4799), .A3(n4238), .A4(n5618), .ZN(n4022)
         );
  BUF_X1 U4055 ( .A(n7104), .Z(n3925) );
  INV_X1 U4056 ( .A(n3925), .ZN(n3926) );
  OR2_X2 U4057 ( .A1(n5176), .A2(\ctrl_u/if_stall ), .ZN(n5626) );
  BUF_X2 U4058 ( .A(n5192), .Z(n3928) );
  OAI21_X1 U4059 ( .B1(n3948), .B2(n4968), .A(n5339), .ZN(n4816) );
  AND2_X2 U4060 ( .A1(n6311), .A2(n6310), .ZN(n6701) );
  INV_X4 U4061 ( .A(n5414), .ZN(n5622) );
  OR2_X2 U4062 ( .A1(n5821), .A2(n6168), .ZN(n5027) );
  AND2_X1 U4063 ( .A1(n4875), .A2(n5044), .ZN(n3931) );
  NAND2_X1 U4064 ( .A1(n4664), .A2(n5023), .ZN(n3932) );
  INV_X1 U4065 ( .A(n3941), .ZN(n3934) );
  BUF_X2 U4066 ( .A(n5192), .Z(n3936) );
  BUF_X2 U4067 ( .A(n7104), .Z(n3937) );
  CLKBUF_X1 U4068 ( .A(n3929), .Z(n4815) );
  BUF_X1 U4069 ( .A(n7439), .Z(n3942) );
  BUF_X2 U4070 ( .A(n7439), .Z(n3938) );
  INV_X1 U4071 ( .A(n7080), .ZN(n3940) );
  AND2_X1 U4072 ( .A1(n5687), .A2(n3899), .ZN(n6298) );
  BUF_X1 U4073 ( .A(n5212), .Z(n3947) );
  NAND2_X2 U4074 ( .A1(n7445), .A2(op_b_fw_sel_exe[0]), .ZN(n7495) );
  OR2_X2 U4075 ( .A1(en_alu_mem), .A2(n5229), .ZN(n7498) );
  INV_X1 U4076 ( .A(n7340), .ZN(n5670) );
  INV_X1 U4077 ( .A(n5156), .ZN(n3944) );
  BUF_X2 U4078 ( .A(n5188), .Z(n3946) );
  BUF_X1 U4079 ( .A(n7083), .Z(n3954) );
  AND2_X2 U4080 ( .A1(n4297), .A2(n5168), .ZN(n6326) );
  NAND2_X1 U4081 ( .A1(n5751), .A2(log_type_exe[3]), .ZN(n7069) );
  BUF_X1 U4082 ( .A(n5212), .Z(n3956) );
  BUF_X1 U4083 ( .A(n7058), .Z(n4048) );
  BUF_X1 U4084 ( .A(n7058), .Z(n4047) );
  BUF_X1 U4085 ( .A(n7179), .Z(n5132) );
  BUF_X1 U4086 ( .A(n7179), .Z(n5131) );
  BUF_X1 U4087 ( .A(n7179), .Z(n5130) );
  NAND2_X1 U4088 ( .A1(n4763), .A2(n4783), .ZN(n4058) );
  NOR2_X1 U4089 ( .A1(n3999), .A2(n4001), .ZN(n3998) );
  BUF_X2 U4090 ( .A(n7491), .Z(n3958) );
  BUF_X2 U4091 ( .A(n7492), .Z(n3959) );
  OAI211_X1 U4092 ( .C1(n6328), .C2(n6103), .A(n6102), .B(n6101), .ZN(n6136)
         );
  OR2_X2 U4093 ( .A1(alu_data_tbs_selector), .A2(n5226), .ZN(n7497) );
  BUF_X1 U4094 ( .A(n7498), .Z(n5227) );
  NOR2_X1 U4095 ( .A1(n5327), .A2(n7251), .ZN(n7064) );
  NAND2_X2 U4096 ( .A1(n4228), .A2(alu_data_tbs_selector), .ZN(n7499) );
  INV_X1 U4097 ( .A(\ctrl_u/n555 ), .ZN(n5339) );
  NOR2_X1 U4098 ( .A1(n5670), .A2(n5229), .ZN(\ctrl_u/n555 ) );
  INV_X2 U4099 ( .A(btb_cache_update_data), .ZN(n6168) );
  NOR2_X1 U4100 ( .A1(n5337), .A2(n5336), .ZN(btb_cache_update_data) );
  INV_X1 U4101 ( .A(n4017), .ZN(n5075) );
  INV_X1 U4102 ( .A(\ctrl_u/mem_stall ), .ZN(n7340) );
  NOR2_X2 U4103 ( .A1(n5686), .A2(n5685), .ZN(n5188) );
  INV_X2 U4104 ( .A(n6157), .ZN(n3952) );
  INV_X1 U4105 ( .A(n7069), .ZN(n3953) );
  NOR2_X4 U4106 ( .A1(n4266), .A2(\mc/currstate[0] ), .ZN(n5191) );
  AND2_X1 U4107 ( .A1(n4297), .A2(n3900), .ZN(n5154) );
  NOR2_X1 U4108 ( .A1(\mc/currstate[1] ), .A2(n4371), .ZN(n4015) );
  AND2_X2 U4109 ( .A1(op_type_exe[1]), .A2(op_type_exe[0]), .ZN(n7076) );
  INV_X1 U4110 ( .A(n5581), .ZN(n5181) );
  OAI21_X1 U4111 ( .B1(n5429), .B2(n4547), .A(n3976), .ZN(\ctrl_u/n521 ) );
  OAI21_X1 U4112 ( .B1(n5429), .B2(n4602), .A(n3976), .ZN(\ctrl_u/n549 ) );
  OAI21_X1 U4113 ( .B1(n5488), .B2(n5560), .A(n5547), .ZN(n5489) );
  BUF_X2 U4114 ( .A(n7057), .Z(n4049) );
  BUF_X2 U4115 ( .A(n7057), .Z(n4050) );
  BUF_X2 U4116 ( .A(n7057), .Z(n4051) );
  INV_X1 U4117 ( .A(n6701), .ZN(n6714) );
  AND2_X1 U4118 ( .A1(n7151), .A2(n4448), .ZN(n4097) );
  OR2_X2 U4119 ( .A1(n7141), .A2(en_imm_id), .ZN(n7163) );
  NAND2_X1 U4120 ( .A1(n4651), .A2(n4933), .ZN(n5653) );
  NOR3_X1 U4121 ( .A1(n7141), .A2(n4396), .A3(n7140), .ZN(n7164) );
  BUF_X1 U4122 ( .A(n7177), .Z(n5133) );
  BUF_X1 U4123 ( .A(n4069), .Z(n5207) );
  INV_X1 U4124 ( .A(n7151), .ZN(n4865) );
  BUF_X1 U4125 ( .A(n7098), .Z(n5126) );
  INV_X2 U4126 ( .A(n6165), .ZN(n5117) );
  BUF_X1 U4127 ( .A(n4107), .Z(n5217) );
  INV_X1 U4128 ( .A(n5215), .ZN(n3955) );
  BUF_X1 U4129 ( .A(n7056), .Z(n5200) );
  BUF_X1 U4130 ( .A(n4069), .Z(n5206) );
  BUF_X1 U4131 ( .A(n7056), .Z(n5201) );
  BUF_X1 U4132 ( .A(n4069), .Z(n5209) );
  BUF_X1 U4133 ( .A(n7177), .Z(n5134) );
  BUF_X1 U4134 ( .A(n4069), .Z(n5210) );
  BUF_X1 U4135 ( .A(n7098), .Z(n5127) );
  BUF_X1 U4136 ( .A(n4069), .Z(n5208) );
  NOR2_X1 U4137 ( .A1(n4820), .A2(n6981), .ZN(n4648) );
  OR2_X1 U4138 ( .A1(n7141), .A2(en_shift_id), .ZN(n7057) );
  BUF_X1 U4139 ( .A(n4107), .Z(n5216) );
  BUF_X1 U4140 ( .A(n5212), .Z(n5211) );
  AND2_X1 U4141 ( .A1(n3901), .A2(n4134), .ZN(n5213) );
  AND2_X2 U4142 ( .A1(n3932), .A2(n4855), .ZN(n4224) );
  AND2_X2 U4143 ( .A1(n3932), .A2(n4316), .ZN(n4107) );
  NAND2_X4 U4144 ( .A1(n3901), .A2(n6334), .ZN(n5199) );
  NOR2_X1 U4145 ( .A1(n5044), .A2(n6171), .ZN(n6165) );
  AND2_X2 U4146 ( .A1(n7171), .A2(n6334), .ZN(n7098) );
  NAND2_X1 U4147 ( .A1(n7005), .A2(n4357), .ZN(n7039) );
  INV_X1 U4148 ( .A(n3873), .ZN(n6405) );
  BUF_X1 U4149 ( .A(n7060), .Z(n5204) );
  OAI21_X1 U4150 ( .B1(n4967), .B2(n3948), .A(n4966), .ZN(n5176) );
  NAND2_X1 U4151 ( .A1(n4816), .A2(pc_en), .ZN(n7179) );
  AND2_X2 U4152 ( .A1(n4965), .A2(n4964), .ZN(n7177) );
  AND2_X1 U4153 ( .A1(n4873), .A2(n4874), .ZN(n6180) );
  OR2_X2 U4154 ( .A1(n6183), .A2(taken), .ZN(n7109) );
  BUF_X1 U4155 ( .A(n7060), .Z(n5203) );
  NAND2_X1 U4156 ( .A1(n3929), .A2(n4922), .ZN(n5416) );
  INV_X2 U4157 ( .A(n5347), .ZN(n5621) );
  BUF_X1 U4158 ( .A(n7060), .Z(n5205) );
  AND2_X1 U4159 ( .A1(n4011), .A2(n4012), .ZN(n4060) );
  OAI21_X1 U4160 ( .B1(n3981), .B2(n7340), .A(n5822), .ZN(n5045) );
  XNOR2_X1 U4161 ( .A(n3967), .B(n3966), .ZN(n4039) );
  NAND2_X1 U4162 ( .A1(\add_x_20/n2 ), .A2(btb_cache_read_address[28]), .ZN(
        n3967) );
  XNOR2_X1 U4163 ( .A(\add_x_20/n2 ), .B(n3869), .ZN(
        \dp/pc_plus4_out_if_int[28] ) );
  CLKBUF_X1 U4164 ( .A(n5052), .Z(n5051) );
  OAI21_X1 U4165 ( .B1(n5923), .B2(n3994), .A(n3993), .ZN(n4782) );
  OAI21_X1 U4166 ( .B1(n5923), .B2(n5089), .A(n4001), .ZN(n4992) );
  OAI21_X1 U4167 ( .B1(n5923), .B2(n5090), .A(n3999), .ZN(n4993) );
  AND3_X1 U4168 ( .A1(\intadd_1/SUM[15] ), .A2(\intadd_1/SUM[8] ), .A3(
        \intadd_1/SUM[9] ), .ZN(n3984) );
  AOI21_X1 U4169 ( .B1(n3995), .B2(n3998), .A(n4058), .ZN(n3993) );
  INV_X1 U4170 ( .A(n3995), .ZN(n3994) );
  INV_X1 U4171 ( .A(\intadd_2/n11 ), .ZN(n3957) );
  AOI21_X1 U4172 ( .B1(n5090), .B2(n3999), .A(n3996), .ZN(n3995) );
  NAND2_X1 U4173 ( .A1(n4951), .A2(n3997), .ZN(n3996) );
  OR2_X1 U4174 ( .A1(n6163), .A2(n4317), .ZN(n5050) );
  NAND2_X1 U4175 ( .A1(n4001), .A2(n5089), .ZN(n3997) );
  NAND2_X2 U4176 ( .A1(n7087), .A2(n7076), .ZN(n7062) );
  NAND2_X2 U4177 ( .A1(n7087), .A2(n5754), .ZN(n7440) );
  OAI21_X1 U4178 ( .B1(n4923), .B2(n3980), .A(n3979), .ZN(\intadd_2/n13 ) );
  XNOR2_X1 U4179 ( .A(n3855), .B(n3867), .ZN(\intadd_2/SUM[15] ) );
  NOR2_X1 U4180 ( .A1(n5333), .A2(n6162), .ZN(n4322) );
  NAND2_X1 U4181 ( .A1(n4751), .A2(\intadd_1/n57 ), .ZN(n4298) );
  OR2_X1 U4182 ( .A1(\intadd_1/A[24] ), .A2(\intadd_1/B[24] ), .ZN(
        \intadd_1/n37 ) );
  OR2_X1 U4183 ( .A1(n5755), .A2(n5229), .ZN(n7439) );
  AND2_X1 U4184 ( .A1(n5755), .A2(rst_mem_wb_regs), .ZN(n7087) );
  OAI21_X1 U4185 ( .B1(n3989), .B2(n3940), .A(n3988), .ZN(n5813) );
  BUF_X1 U4186 ( .A(n7108), .Z(n5193) );
  BUF_X1 U4187 ( .A(en_shift_id), .Z(n6473) );
  INV_X1 U4188 ( .A(n5024), .ZN(n5023) );
  INV_X1 U4189 ( .A(n7391), .ZN(n7394) );
  NAND2_X1 U4190 ( .A1(n3989), .A2(n7069), .ZN(n3988) );
  NOR3_X1 U4191 ( .A1(n5925), .A2(n5092), .A3(n5089), .ZN(n4994) );
  OAI211_X1 U4192 ( .C1(n6328), .C2(n6093), .A(n6092), .B(n6091), .ZN(n6099)
         );
  NOR2_X1 U4193 ( .A1(n5026), .A2(n5339), .ZN(n5024) );
  OAI21_X1 U4194 ( .B1(n7260), .B2(n4264), .A(n7259), .ZN(n92) );
  INV_X1 U4195 ( .A(n6333), .ZN(n5026) );
  AND2_X1 U4196 ( .A1(n7397), .A2(n7396), .ZN(n7413) );
  INV_X1 U4197 ( .A(n7381), .ZN(n7383) );
  INV_X1 U4198 ( .A(n7414), .ZN(n7392) );
  NAND2_X1 U4199 ( .A1(n5421), .A2(n5420), .ZN(\ctrl_u/if_stall ) );
  AND2_X1 U4200 ( .A1(n7298), .A2(\ctrl_u/curr_exe[16] ), .ZN(en_b_exe) );
  NOR2_X1 U4201 ( .A1(n7382), .A2(n7381), .ZN(n7396) );
  OAI211_X1 U4202 ( .C1(n3930), .C2(n4064), .A(n6095), .B(n6094), .ZN(n6100)
         );
  AND2_X1 U4203 ( .A1(rst_mem_wb_regs), .A2(en_alu_mem), .ZN(n4228) );
  NOR2_X1 U4204 ( .A1(n5769), .A2(n4300), .ZN(op_b_fw_sel_exe[0]) );
  OR2_X1 U4205 ( .A1(n5669), .A2(n5668), .ZN(n7338) );
  BUF_X1 U4206 ( .A(n7253), .Z(n5174) );
  INV_X1 U4207 ( .A(n5822), .ZN(n5824) );
  BUF_X1 U4208 ( .A(n5140), .Z(n4043) );
  BUF_X1 U4209 ( .A(n5136), .Z(n4016) );
  AND2_X1 U4210 ( .A1(n5655), .A2(n5670), .ZN(n5420) );
  AND2_X1 U4211 ( .A1(n5670), .A2(\ctrl_u/curr_mem[6] ), .ZN(en_alu_mem) );
  AND2_X1 U4212 ( .A1(n5670), .A2(\ctrl_u/curr_mem[5] ), .ZN(en_cache_mem) );
  INV_X1 U4213 ( .A(n5655), .ZN(n5413) );
  NOR2_X2 U4214 ( .A1(n5620), .A2(\ctrl_u/curr_mul_in_prog ), .ZN(n5655) );
  INV_X1 U4215 ( .A(n6323), .ZN(n3960) );
  BUF_X1 U4216 ( .A(n5098), .Z(n4037) );
  AOI21_X1 U4217 ( .B1(n5232), .B2(\ctrl_u/curr_ms ), .A(n5231), .ZN(
        \ctrl_u/mem_stall ) );
  AND2_X1 U4218 ( .A1(n5054), .A2(n5078), .ZN(n4017) );
  NOR2_X1 U4219 ( .A1(n6327), .A2(n7274), .ZN(n5753) );
  INV_X2 U4220 ( .A(n3113), .ZN(n7425) );
  INV_X1 U4221 ( .A(n5086), .ZN(n3961) );
  BUF_X2 U4222 ( .A(n5183), .Z(n3963) );
  NAND2_X1 U4223 ( .A1(n7188), .A2(n3910), .ZN(n5232) );
  AND4_X1 U4224 ( .A1(n5361), .A2(n5360), .A3(n5359), .A4(n5358), .ZN(n4299)
         );
  INV_X1 U4225 ( .A(n6298), .ZN(n6328) );
  INV_X1 U4226 ( .A(n5061), .ZN(n5231) );
  INV_X1 U4227 ( .A(n3900), .ZN(n6327) );
  INV_X1 U4228 ( .A(n7076), .ZN(n6027) );
  OR2_X1 U4229 ( .A1(n5164), .A2(n5162), .ZN(n5679) );
  INV_X1 U4230 ( .A(n5671), .ZN(n5097) );
  AND2_X1 U4231 ( .A1(n5263), .A2(n5265), .ZN(n3968) );
  OR2_X1 U4232 ( .A1(n4015), .A2(n5088), .ZN(n4740) );
  XNOR2_X1 U4233 ( .A(\add_x_20/n28 ), .B(n3868), .ZN(
        \dp/pc_plus4_out_if_int[2] ) );
  AND2_X1 U4234 ( .A1(\add_x_20/n28 ), .A2(btb_cache_read_address[2]), .ZN(
        \add_x_20/n27 ) );
  NOR2_X2 U4235 ( .A1(n4266), .A2(\mc/currstate[0] ), .ZN(n5810) );
  NAND2_X1 U4236 ( .A1(n4257), .A2(n4113), .ZN(n3979) );
  AND2_X1 U4237 ( .A1(cpu_is_reading), .A2(n4127), .ZN(n5063) );
  NOR2_X1 U4238 ( .A1(n4257), .A2(n4113), .ZN(n3980) );
  INV_X1 U4239 ( .A(n5161), .ZN(n5162) );
  INV_X1 U4240 ( .A(n5163), .ZN(n5164) );
  CLKBUF_X1 U4241 ( .A(rd_exemem[1]), .Z(n3970) );
  INV_X1 U4242 ( .A(n4005), .ZN(rd[1]) );
  CLKBUF_X1 U4243 ( .A(n7535), .Z(rd[3]) );
  BUF_X1 U4244 ( .A(n7536), .Z(rd[2]) );
  BUF_X1 U4245 ( .A(n7534), .Z(rd[4]) );
  BUF_X1 U4246 ( .A(n7538), .Z(rd[0]) );
  INV_X1 U4247 ( .A(n4358), .ZN(n5230) );
  NOR2_X1 U4248 ( .A1(op_type_exe[1]), .A2(op_type_exe[0]), .ZN(n7083) );
  INV_X1 U4249 ( .A(n5552), .ZN(n3962) );
  INV_X1 U4250 ( .A(instr_if[1]), .ZN(n7280) );
  INV_X1 U4251 ( .A(cache_to_ram_data[19]), .ZN(n7510) );
  INV_X1 U4252 ( .A(cache_to_ram_data[28]), .ZN(n7520) );
  INV_X1 U4253 ( .A(instr_if[29]), .ZN(n7275) );
  INV_X1 U4254 ( .A(cache_to_ram_data[20]), .ZN(n7512) );
  INV_X1 U4255 ( .A(cache_to_ram_data[26]), .ZN(n7518) );
  INV_X1 U4256 ( .A(instr_if[0]), .ZN(n7281) );
  INV_X1 U4257 ( .A(cache_to_ram_data[25]), .ZN(n7517) );
  INV_X1 U4258 ( .A(cache_to_ram_data[21]), .ZN(n7513) );
  INV_X1 U4259 ( .A(instr_if[2]), .ZN(n5530) );
  INV_X1 U4260 ( .A(instr_if[5]), .ZN(n7277) );
  INV_X1 U4261 ( .A(cache_to_ram_data[23]), .ZN(n7515) );
  INV_X1 U4262 ( .A(cache_to_ram_data[22]), .ZN(n7514) );
  INV_X1 U4263 ( .A(cache_to_ram_data[24]), .ZN(n7516) );
  INV_X1 U4264 ( .A(cache_to_ram_data[27]), .ZN(n7519) );
  INV_X1 U4265 ( .A(cache_to_ram_data[30]), .ZN(n7523) );
  INV_X1 U4266 ( .A(instr_if[31]), .ZN(n5644) );
  INV_X1 U4267 ( .A(cache_to_ram_data[1]), .ZN(n7511) );
  INV_X1 U4268 ( .A(cache_to_ram_data[2]), .ZN(n7522) );
  INV_X1 U4269 ( .A(instr_if[27]), .ZN(n5627) );
  INV_X1 U4270 ( .A(cache_to_ram_data[13]), .ZN(n7504) );
  INV_X1 U4271 ( .A(cache_to_ram_data[3]), .ZN(n7525) );
  INV_X1 U4272 ( .A(instr_if[30]), .ZN(n5590) );
  INV_X1 U4273 ( .A(cache_to_ram_data[4]), .ZN(n7526) );
  INV_X1 U4274 ( .A(cache_to_ram_data[5]), .ZN(n7527) );
  INV_X1 U4275 ( .A(rst_mem_wb_regs), .ZN(n5229) );
  INV_X1 U4276 ( .A(cache_to_ram_data[12]), .ZN(n7503) );
  INV_X1 U4277 ( .A(cache_to_ram_data[6]), .ZN(n7528) );
  INV_X1 U4278 ( .A(cache_to_ram_data[31]), .ZN(n7524) );
  INV_X1 U4279 ( .A(cache_to_ram_data[7]), .ZN(n7529) );
  INV_X1 U4280 ( .A(instr_if[26]), .ZN(n5560) );
  INV_X1 U4281 ( .A(cache_to_ram_data[11]), .ZN(n7502) );
  INV_X1 U4282 ( .A(ram_update), .ZN(n5677) );
  INV_X1 U4283 ( .A(cache_to_ram_data[8]), .ZN(n7530) );
  INV_X1 U4284 ( .A(cache_to_ram_data[10]), .ZN(n7501) );
  INV_X1 U4285 ( .A(cache_to_ram_data[9]), .ZN(n7531) );
  INV_X1 U4286 ( .A(cache_to_ram_data[18]), .ZN(n7509) );
  INV_X1 U4287 ( .A(instr_if[3]), .ZN(n7279) );
  INV_X1 U4288 ( .A(cache_to_ram_data[17]), .ZN(n7508) );
  INV_X1 U4289 ( .A(cache_to_ram_data[29]), .ZN(n7521) );
  INV_X1 U4290 ( .A(cache_to_ram_data[16]), .ZN(n7507) );
  INV_X1 U4291 ( .A(cache_to_ram_data[15]), .ZN(n7506) );
  INV_X1 U4292 ( .A(cache_to_ram_data[0]), .ZN(n7500) );
  INV_X1 U4293 ( .A(cache_to_ram_data[14]), .ZN(n7505) );
  AND2_X1 U4294 ( .A1(btb_addr_known_if), .A2(btb_cache_data_out_read[31]), 
        .ZN(predicted_taken) );
  OAI211_X4 U4295 ( .C1(n5676), .C2(n5675), .A(n5674), .B(n5673), .ZN(n7337)
         );
  NAND2_X1 U4296 ( .A1(n5062), .A2(n3964), .ZN(n5098) );
  NAND2_X1 U4297 ( .A1(n3965), .A2(n3910), .ZN(n3964) );
  INV_X1 U4298 ( .A(n5088), .ZN(n3965) );
  NAND2_X1 U4299 ( .A1(n4703), .A2(n4704), .ZN(n5062) );
  INV_X1 U4300 ( .A(n7171), .ZN(n7141) );
  NAND3_X1 U4301 ( .A1(n4033), .A2(n4859), .A3(n4034), .ZN(n6055) );
  NAND3_X1 U4302 ( .A1(n4836), .A2(n5266), .A3(n3968), .ZN(n5340) );
  NAND2_X2 U4303 ( .A1(n5137), .A2(n3961), .ZN(n5172) );
  NAND2_X1 U4304 ( .A1(n5088), .A2(n5063), .ZN(n5061) );
  NAND3_X1 U4305 ( .A1(n5160), .A2(\ctrl_u/curr_mul_end_wb ), .A3(n5157), .ZN(
        n4762) );
  NAND2_X1 U4306 ( .A1(n5626), .A2(n3929), .ZN(n5652) );
  NAND2_X1 U4307 ( .A1(n3974), .A2(n6403), .ZN(n4661) );
  AOI21_X1 U4308 ( .B1(n3926), .B2(n4662), .A(n3975), .ZN(n3974) );
  NOR2_X1 U4309 ( .A1(n7109), .A2(n4536), .ZN(n3975) );
  OAI21_X1 U4310 ( .B1(n5429), .B2(n4586), .A(n3976), .ZN(\ctrl_u/n542 ) );
  NAND2_X1 U4311 ( .A1(n3978), .A2(n3977), .ZN(n3976) );
  NOR2_X1 U4312 ( .A1(\ctrl_u/if_stall ), .A2(n5428), .ZN(n3977) );
  INV_X1 U4313 ( .A(n5130), .ZN(n3978) );
  NAND2_X1 U4314 ( .A1(n7533), .A2(\ctrl_u/curr_exe_41 ), .ZN(n3981) );
  NAND2_X1 U4315 ( .A1(n3982), .A2(n4721), .ZN(n7533) );
  OAI21_X1 U4316 ( .B1(n4879), .B2(n4723), .A(n4722), .ZN(n3982) );
  NOR2_X1 U4317 ( .A1(n3985), .A2(n3983), .ZN(n4769) );
  NAND4_X1 U4318 ( .A1(\intadd_1/SUM[14] ), .A2(n3984), .A3(\intadd_1/SUM[25] ), .A4(\intadd_1/SUM[19] ), .ZN(n3983) );
  NAND2_X1 U4319 ( .A1(\intadd_1/SUM[18] ), .A2(\intadd_1/SUM[26] ), .ZN(n3985) );
  XNOR2_X1 U4320 ( .A(n3986), .B(n4777), .ZN(\intadd_1/SUM[26] ) );
  OAI21_X1 U4321 ( .B1(n4725), .B2(n4724), .A(n5076), .ZN(n3986) );
  XNOR2_X1 U4322 ( .A(n3987), .B(\intadd_1/n8 ), .ZN(\intadd_1/SUM[18] ) );
  OAI21_X1 U4323 ( .B1(n4761), .B2(n3860), .A(\intadd_1/n78 ), .ZN(n3987) );
  XNOR2_X1 U4324 ( .A(n3989), .B(sub_add_exe), .ZN(\intadd_1/B[1] ) );
  NAND2_X1 U4325 ( .A1(n5323), .A2(n7257), .ZN(n3989) );
  OR2_X1 U4326 ( .A1(n5140), .A2(n3990), .ZN(n3991) );
  OR2_X1 U4327 ( .A1(n5141), .A2(\dp/b_adder_id_exe_int[11] ), .ZN(n3990) );
  AND2_X1 U4328 ( .A1(n5253), .A2(n3991), .ZN(n5109) );
  XNOR2_X1 U4329 ( .A(n3992), .B(n4225), .ZN(\intadd_1/A[9] ) );
  NAND2_X1 U4330 ( .A1(n5255), .A2(n5254), .ZN(n3992) );
  NOR2_X1 U4331 ( .A1(n4994), .A2(n4000), .ZN(n3999) );
  INV_X1 U4332 ( .A(n5926), .ZN(n4000) );
  INV_X1 U4333 ( .A(n4003), .ZN(n4004) );
  OAI22_X1 U4334 ( .A1(n4039), .A2(n7105), .B1(n3873), .B2(n4483), .ZN(n4003)
         );
  INV_X1 U4335 ( .A(n4007), .ZN(n4008) );
  INV_X1 U4336 ( .A(n4009), .ZN(n4010) );
  NAND2_X1 U4337 ( .A1(n6088), .A2(n4014), .ZN(n4011) );
  OR2_X1 U4338 ( .A1(n4013), .A2(n4716), .ZN(n4012) );
  INV_X1 U4339 ( .A(n6100), .ZN(n4013) );
  AND2_X1 U4340 ( .A1(n4309), .A2(n6100), .ZN(n4014) );
  NOR2_X1 U4341 ( .A1(\intadd_1/A[12] ), .A2(\intadd_1/B[12] ), .ZN(
        \intadd_1/n109 ) );
  AND4_X1 U4342 ( .A1(n4960), .A2(n4841), .A3(\ctrl_u/curr_mem[3] ), .A4(n5239), .ZN(n4728) );
  CLKBUF_X1 U4343 ( .A(n7533), .Z(taken) );
  INV_X1 U4344 ( .A(n4018), .ZN(n4019) );
  INV_X1 U4345 ( .A(n4020), .ZN(n4021) );
  NOR2_X1 U4346 ( .A1(n3910), .A2(n5678), .ZN(n3113) );
  OAI21_X1 U4347 ( .B1(n3910), .B2(n5677), .A(rst_mem_wb_regs), .ZN(n5183) );
  INV_X1 U4348 ( .A(n7179), .ZN(n7186) );
  AOI21_X1 U4349 ( .B1(n4872), .B2(n5027), .A(n4328), .ZN(n7060) );
  NOR2_X1 U4350 ( .A1(n7141), .A2(en_rd_id), .ZN(n7166) );
  OR4_X1 U4351 ( .A1(n5653), .A2(n5548), .A3(n3962), .A4(instr_if[27]), .ZN(
        n5554) );
  NAND3_X1 U4352 ( .A1(n3907), .A2(n4060), .A3(n4061), .ZN(n4023) );
  NAND3_X1 U4353 ( .A1(n4059), .A2(n4060), .A3(n4061), .ZN(n6148) );
  INV_X1 U4354 ( .A(n5160), .ZN(n4025) );
  NOR2_X1 U4355 ( .A1(\intadd_1/B[20] ), .A2(n4845), .ZN(n4026) );
  AOI21_X1 U4356 ( .B1(n5135), .B2(n4304), .A(n4702), .ZN(n6012) );
  INV_X1 U4357 ( .A(n5626), .ZN(n5599) );
  INV_X1 U4358 ( .A(n5170), .ZN(n7260) );
  INV_X1 U4359 ( .A(n4832), .ZN(n4027) );
  AND2_X1 U4360 ( .A1(n3884), .A2(n6410), .ZN(n4028) );
  OAI21_X1 U4361 ( .B1(\intadd_1/n171 ), .B2(\intadd_1/n173 ), .A(
        \intadd_1/n172 ), .ZN(n4029) );
  XNOR2_X1 U4362 ( .A(n4725), .B(n4030), .ZN(\intadd_1/SUM[24] ) );
  AND2_X1 U4363 ( .A1(\intadd_1/n37 ), .A2(\intadd_1/n38 ), .ZN(n4030) );
  BUF_X1 U4364 ( .A(n5768), .Z(n4031) );
  BUF_X1 U4365 ( .A(n3922), .Z(n4041) );
  AND2_X1 U4366 ( .A1(\ctrl_u/n95 ), .A2(\ctrl_u/n94 ), .ZN(n7273) );
  INV_X1 U4367 ( .A(n3957), .ZN(n4032) );
  NAND2_X1 U4368 ( .A1(n5969), .A2(n4036), .ZN(n4033) );
  OR2_X1 U4369 ( .A1(n4035), .A2(n4800), .ZN(n4034) );
  INV_X1 U4370 ( .A(n4857), .ZN(n4035) );
  AND2_X1 U4371 ( .A1(n4310), .A2(n4857), .ZN(n4036) );
  NAND2_X1 U4372 ( .A1(n4874), .A2(n6176), .ZN(n5044) );
  XNOR2_X1 U4373 ( .A(n5109), .B(sub_add_exe), .ZN(n4038) );
  AOI21_X1 U4374 ( .B1(n4720), .B2(\intadd_1/n120 ), .A(\intadd_1/n121 ), .ZN(
        \intadd_1/n119 ) );
  INV_X1 U4375 ( .A(n5140), .ZN(n5273) );
  BUF_X1 U4376 ( .A(n5882), .Z(n4042) );
  XNOR2_X1 U4377 ( .A(n6527), .B(n4044), .ZN(n6528) );
  AND2_X1 U4378 ( .A1(n6519), .A2(n6518), .ZN(n4044) );
  OR2_X1 U4379 ( .A1(\intadd_1/A[2] ), .A2(\intadd_1/B[2] ), .ZN(n4045) );
  XNOR2_X1 U4380 ( .A(n6539), .B(n4046), .ZN(n6540) );
  AND2_X1 U4381 ( .A1(n6533), .A2(n6532), .ZN(n4046) );
  XNOR2_X1 U4382 ( .A(n6603), .B(n4053), .ZN(n6604) );
  AND2_X1 U4383 ( .A1(n6598), .A2(n6597), .ZN(n4053) );
  NAND2_X1 U4384 ( .A1(n3933), .A2(\ctrl_u/n83 ), .ZN(n5336) );
  AND2_X1 U4385 ( .A1(n5157), .A2(n4025), .ZN(n7274) );
  INV_X1 U4386 ( .A(n5157), .ZN(n5158) );
  NAND2_X1 U4387 ( .A1(n4799), .A2(n5234), .ZN(n5620) );
  NAND2_X1 U4388 ( .A1(n6098), .A2(n6099), .ZN(n4059) );
  NAND2_X1 U4389 ( .A1(n6099), .A2(n6100), .ZN(n4061) );
  NAND2_X1 U4390 ( .A1(n4871), .A2(n5027), .ZN(n4664) );
  NOR2_X1 U4391 ( .A1(n4266), .A2(\mc/currstate[0] ), .ZN(n5190) );
  OR2_X1 U4392 ( .A1(n3927), .A2(n4604), .ZN(n5571) );
  OR2_X1 U4393 ( .A1(n3927), .A2(n4856), .ZN(n5570) );
  INV_X1 U4394 ( .A(n5653), .ZN(n5641) );
  NOR2_X1 U4395 ( .A1(\intadd_1/n127 ), .A2(n4706), .ZN(\intadd_1/n120 ) );
  AND2_X1 U4396 ( .A1(n3932), .A2(n4843), .ZN(n4069) );
  AND2_X1 U4397 ( .A1(n7171), .A2(n4353), .ZN(n5212) );
  NOR2_X4 U4398 ( .A1(en_cache_mem), .A2(n5229), .ZN(n7414) );
  AOI21_X2 U4399 ( .B1(ld_sign_mem), .B2(n7395), .A(n7394), .ZN(n7416) );
  NOR2_X4 U4400 ( .A1(op_b_fw_sel_exe[0]), .A2(n7446), .ZN(n7493) );
  OAI21_X1 U4401 ( .B1(n7150), .B2(n7148), .A(n7151), .ZN(n7149) );
  BUF_X2 U4402 ( .A(n7163), .Z(n5224) );
  NAND2_X1 U4403 ( .A1(n7151), .A2(n7150), .ZN(n7161) );
  BUF_X2 U4404 ( .A(n7163), .Z(n5225) );
  INV_X1 U4405 ( .A(n5195), .ZN(n5197) );
  BUF_X1 U4406 ( .A(n7139), .Z(n5218) );
  BUF_X1 U4407 ( .A(n7139), .Z(n5222) );
  BUF_X1 U4408 ( .A(n7139), .Z(n5219) );
  BUF_X1 U4409 ( .A(n7139), .Z(n5221) );
  BUF_X1 U4410 ( .A(n7139), .Z(n5220) );
  BUF_X1 U4411 ( .A(n7139), .Z(n5223) );
  INV_X1 U4412 ( .A(n5549), .ZN(n5565) );
  AND2_X1 U4413 ( .A1(n6310), .A2(n6311), .ZN(n5125) );
  NAND2_X1 U4414 ( .A1(n4850), .A2(n4844), .ZN(n5563) );
  INV_X1 U4415 ( .A(n5195), .ZN(n5198) );
  INV_X1 U4416 ( .A(n6719), .ZN(n5195) );
  BUF_X1 U4417 ( .A(n7056), .Z(n5202) );
  NAND2_X1 U4418 ( .A1(n7097), .A2(n7076), .ZN(n6719) );
  NAND2_X1 U4419 ( .A1(n6309), .A2(n6308), .ZN(n6310) );
  AOI21_X1 U4420 ( .B1(n6148), .B2(n6147), .A(n6146), .ZN(n6309) );
  NOR2_X1 U4421 ( .A1(n7060), .A2(n6981), .ZN(n6991) );
  NOR2_X1 U4422 ( .A1(n7060), .A2(n4357), .ZN(n7036) );
  AND2_X1 U4423 ( .A1(n4968), .A2(n5339), .ZN(n4821) );
  AOI21_X1 U4424 ( .B1(n4868), .B2(n5027), .A(n4866), .ZN(n5347) );
  NAND2_X1 U4425 ( .A1(n4717), .A2(n4716), .ZN(n6098) );
  NAND2_X2 U4426 ( .A1(n4236), .A2(op_type_exe[1]), .ZN(n7066) );
  OR2_X1 U4427 ( .A1(n6029), .A2(n6030), .ZN(n5077) );
  NAND2_X1 U4428 ( .A1(n4801), .A2(n4800), .ZN(n5988) );
  AND2_X1 U4429 ( .A1(n5757), .A2(n5756), .ZN(n4106) );
  AND2_X1 U4430 ( .A1(n5725), .A2(n5726), .ZN(n5888) );
  OR2_X1 U4431 ( .A1(n5149), .A2(n5155), .ZN(n5680) );
  INV_X1 U4432 ( .A(n6183), .ZN(n6179) );
  OR2_X1 U4433 ( .A1(n6176), .A2(n6181), .ZN(n6183) );
  NAND3_X1 U4434 ( .A1(n5046), .A2(n5823), .A3(n5045), .ZN(n6176) );
  BUF_X2 U4435 ( .A(n5213), .Z(n5214) );
  NAND2_X1 U4436 ( .A1(n6923), .A2(n6980), .ZN(n6958) );
  INV_X1 U4437 ( .A(n6931), .ZN(n7100) );
  INV_X1 U4438 ( .A(n7177), .ZN(n5178) );
  AOI21_X1 U4439 ( .B1(n3858), .B2(n5339), .A(pc_en), .ZN(n4964) );
  OAI21_X1 U4440 ( .B1(n4854), .B2(n3948), .A(n4117), .ZN(n4933) );
  OR2_X1 U4441 ( .A1(n4968), .A2(pc_en), .ZN(n4967) );
  XNOR2_X1 U4442 ( .A(n7533), .B(\ctrl_u/curr_pt_exe ), .ZN(n5821) );
  AND2_X1 U4443 ( .A1(n5338), .A2(n5025), .ZN(n4871) );
  OAI211_X1 U4444 ( .C1(n5143), .C2(n4126), .A(n4944), .B(n4349), .ZN(n4721)
         );
  OR2_X1 U4445 ( .A1(n7092), .A2(n4126), .ZN(n4349) );
  AOI21_X1 U4446 ( .B1(n7092), .B2(n4126), .A(cond_sel_exe[2]), .ZN(n4944) );
  OAI21_X1 U4447 ( .B1(n5143), .B2(n4945), .A(n4494), .ZN(n4722) );
  NAND2_X1 U4448 ( .A1(n4989), .A2(n4771), .ZN(n5143) );
  AND2_X1 U4449 ( .A1(n4906), .A2(n4981), .ZN(n4771) );
  AND2_X1 U4450 ( .A1(n5052), .A2(n5043), .ZN(n4723) );
  OAI21_X1 U4451 ( .B1(cond_sel_exe[0]), .B2(n5052), .A(n5042), .ZN(n4879) );
  NAND2_X1 U4452 ( .A1(n4989), .A2(n4766), .ZN(n5052) );
  AND2_X1 U4453 ( .A1(\intadd_1/SUM[22] ), .A2(n4790), .ZN(n4764) );
  AND2_X1 U4454 ( .A1(\intadd_1/SUM[12] ), .A2(\intadd_1/SUM[20] ), .ZN(n4790)
         );
  OAI21_X1 U4455 ( .B1(n4760), .B2(n4754), .A(n4752), .ZN(\intadd_1/n55 ) );
  AND2_X1 U4456 ( .A1(n4301), .A2(\intadd_1/SUM[28] ), .ZN(n4765) );
  OAI211_X1 U4457 ( .C1(n4789), .C2(n4708), .A(n4707), .B(n4331), .ZN(
        \intadd_1/SUM[28] ) );
  AND4_X1 U4458 ( .A1(\intadd_1/SUM[17] ), .A2(\intadd_1/SUM[13] ), .A3(
        \intadd_1/SUM[23] ), .A4(\intadd_1/SUM[16] ), .ZN(n4301) );
  AOI21_X1 U4459 ( .B1(\intadd_1/n89 ), .B2(\intadd_1/n80 ), .A(\intadd_1/n81 ), .ZN(n4761) );
  OAI21_X1 U4460 ( .B1(\intadd_1/n139 ), .B2(n4833), .A(n4831), .ZN(
        \intadd_1/n104 ) );
  NOR2_X1 U4461 ( .A1(n4768), .A2(n4770), .ZN(n4767) );
  INV_X1 U4462 ( .A(\intadd_1/n69 ), .ZN(n5060) );
  INV_X1 U4463 ( .A(\intadd_1/n71 ), .ZN(\intadd_1/n69 ) );
  INV_X1 U4464 ( .A(\intadd_1/n70 ), .ZN(\intadd_1/n68 ) );
  INV_X1 U4465 ( .A(\intadd_1/n89 ), .ZN(n4760) );
  INV_X1 U4466 ( .A(\intadd_1/n90 ), .ZN(\intadd_1/n89 ) );
  NAND4_X1 U4467 ( .A1(n4791), .A2(\intadd_1/SUM[10] ), .A3(n4128), .A4(
        \intadd_1/SUM[6] ), .ZN(n4768) );
  AND4_X1 U4468 ( .A1(n4302), .A2(\intadd_1/SUM[7] ), .A3(\intadd_1/SUM[5] ), 
        .A4(n4995), .ZN(n4128) );
  AND3_X1 U4469 ( .A1(n5329), .A2(\intadd_1/SUM[3] ), .A3(\intadd_1/SUM[2] ), 
        .ZN(n4302) );
  OAI21_X1 U4470 ( .B1(\intadd_1/n139 ), .B2(\intadd_1/n130 ), .A(
        \intadd_1/n131 ), .ZN(n4729) );
  AND2_X1 U4471 ( .A1(\intadd_1/SUM[24] ), .A2(\intadd_1/SUM[11] ), .ZN(n4791)
         );
  INV_X1 U4472 ( .A(\intadd_1/n140 ), .ZN(\intadd_1/n139 ) );
  AND2_X1 U4473 ( .A1(\intadd_1/SUM[29] ), .A2(n6164), .ZN(n4766) );
  NOR2_X1 U4474 ( .A1(\intadd_1/A[29] ), .A2(\intadd_1/B[29] ), .ZN(n5070) );
  AND2_X1 U4475 ( .A1(\intadd_1/A[29] ), .A2(\intadd_1/B[29] ), .ZN(n4287) );
  XNOR2_X1 U4476 ( .A(n5333), .B(n6162), .ZN(n5332) );
  NOR2_X1 U4477 ( .A1(n5331), .A2(n7189), .ZN(n6162) );
  NOR2_X1 U4478 ( .A1(n5175), .A2(n494), .ZN(n5331) );
  NOR2_X1 U4479 ( .A1(n5277), .A2(n7191), .ZN(\intadd_1/B[29] ) );
  NAND2_X1 U4480 ( .A1(n5276), .A2(n5275), .ZN(n7191) );
  OR2_X1 U4481 ( .A1(n5172), .A2(n5274), .ZN(n5275) );
  XNOR2_X1 U4482 ( .A(n6124), .B(n4225), .ZN(\intadd_1/A[29] ) );
  INV_X1 U4483 ( .A(n4803), .ZN(n4795) );
  OR2_X1 U4484 ( .A1(\intadd_1/A[27] ), .A2(\intadd_1/B[27] ), .ZN(n4803) );
  NOR2_X1 U4485 ( .A1(n4796), .A2(n4256), .ZN(n4731) );
  AND2_X1 U4486 ( .A1(\intadd_1/A[28] ), .A2(\intadd_1/B[28] ), .ZN(n4256) );
  NOR2_X1 U4487 ( .A1(n5281), .A2(n7193), .ZN(\intadd_1/B[28] ) );
  XNOR2_X1 U4488 ( .A(n6113), .B(n4225), .ZN(\intadd_1/A[28] ) );
  INV_X1 U4489 ( .A(n4802), .ZN(n4796) );
  NAND2_X1 U4490 ( .A1(\intadd_1/A[27] ), .A2(\intadd_1/B[27] ), .ZN(n4802) );
  NOR2_X1 U4491 ( .A1(n5283), .A2(n7195), .ZN(\intadd_1/B[27] ) );
  XNOR2_X1 U4492 ( .A(n6105), .B(n4225), .ZN(\intadd_1/A[27] ) );
  NAND2_X1 U4493 ( .A1(\intadd_1/n33 ), .A2(n4700), .ZN(n4709) );
  NAND2_X1 U4494 ( .A1(\intadd_1/n36 ), .A2(n4229), .ZN(n4700) );
  INV_X1 U4495 ( .A(\intadd_1/n38 ), .ZN(\intadd_1/n36 ) );
  NAND3_X1 U4496 ( .A1(n4352), .A2(n4229), .A3(\intadd_1/n39 ), .ZN(n4732) );
  OAI21_X1 U4497 ( .B1(\intadd_1/n90 ), .B2(\intadd_1/n40 ), .A(\intadd_1/n41 ), .ZN(\intadd_1/n39 ) );
  AOI21_X1 U4498 ( .B1(\intadd_1/n48 ), .B2(n4208), .A(\intadd_1/n43 ), .ZN(
        \intadd_1/n41 ) );
  OAI21_X1 U4499 ( .B1(\intadd_1/n49 ), .B2(\intadd_1/n71 ), .A(\intadd_1/n50 ), .ZN(\intadd_1/n48 ) );
  AOI21_X1 U4500 ( .B1(\intadd_1/n72 ), .B2(\intadd_1/n81 ), .A(\intadd_1/n73 ), .ZN(\intadd_1/n71 ) );
  NAND2_X1 U4501 ( .A1(\intadd_1/n47 ), .A2(n4208), .ZN(\intadd_1/n40 ) );
  OR2_X1 U4502 ( .A1(\intadd_1/A[23] ), .A2(\intadd_1/B[23] ), .ZN(n4208) );
  XNOR2_X1 U4503 ( .A(n6047), .B(sub_add_exe), .ZN(\intadd_1/A[23] ) );
  AOI21_X1 U4504 ( .B1(n5170), .B2(n4342), .A(n5241), .ZN(n6047) );
  NOR2_X1 U4505 ( .A1(\intadd_1/n49 ), .A2(\intadd_1/n70 ), .ZN(\intadd_1/n47 ) );
  NAND2_X1 U4506 ( .A1(\intadd_1/n80 ), .A2(\intadd_1/n72 ), .ZN(
        \intadd_1/n70 ) );
  NOR2_X1 U4507 ( .A1(\intadd_1/n77 ), .A2(\intadd_1/n74 ), .ZN(\intadd_1/n72 ) );
  AOI21_X1 U4508 ( .B1(n5118), .B2(n4248), .A(n7213), .ZN(\intadd_1/B[18] ) );
  XNOR2_X1 U4509 ( .A(n5978), .B(sub_add_exe), .ZN(\intadd_1/A[18] ) );
  AOI21_X1 U4510 ( .B1(n5122), .B2(n4339), .A(n5244), .ZN(n5978) );
  NOR2_X1 U4511 ( .A1(\intadd_1/A[17] ), .A2(\intadd_1/B[17] ), .ZN(
        \intadd_1/n77 ) );
  AOI21_X1 U4512 ( .B1(n5118), .B2(n4249), .A(n7215), .ZN(\intadd_1/B[17] ) );
  AOI21_X1 U4513 ( .B1(n5122), .B2(n4338), .A(n5245), .ZN(n5961) );
  NOR2_X1 U4514 ( .A1(\intadd_1/n87 ), .A2(\intadd_1/n82 ), .ZN(\intadd_1/n80 ) );
  NOR2_X1 U4515 ( .A1(\intadd_1/A[16] ), .A2(\intadd_1/B[16] ), .ZN(
        \intadd_1/n82 ) );
  NOR2_X1 U4516 ( .A1(n5298), .A2(n7217), .ZN(\intadd_1/B[16] ) );
  XNOR2_X1 U4517 ( .A(n5760), .B(n4225), .ZN(\intadd_1/A[16] ) );
  NAND2_X1 U4518 ( .A1(n5247), .A2(n5246), .ZN(n5760) );
  NOR2_X1 U4519 ( .A1(n5300), .A2(n7219), .ZN(\intadd_1/B[15] ) );
  NAND2_X1 U4520 ( .A1(\intadd_1/n59 ), .A2(\intadd_1/n51 ), .ZN(
        \intadd_1/n49 ) );
  NOR2_X1 U4521 ( .A1(\intadd_1/n56 ), .A2(\intadd_1/n53 ), .ZN(\intadd_1/n51 ) );
  NOR2_X1 U4522 ( .A1(n4699), .A2(\intadd_1/B[22] ), .ZN(\intadd_1/n53 ) );
  NOR2_X1 U4523 ( .A1(\intadd_1/A[21] ), .A2(\intadd_1/B[21] ), .ZN(
        \intadd_1/n56 ) );
  AOI21_X1 U4524 ( .B1(n5118), .B2(n4245), .A(n7207), .ZN(\intadd_1/B[21] ) );
  AND2_X1 U4525 ( .A1(n5120), .A2(n4335), .ZN(n4730) );
  NOR2_X1 U4526 ( .A1(n4845), .A2(\intadd_1/B[20] ), .ZN(\intadd_1/n61 ) );
  NOR2_X1 U4527 ( .A1(\intadd_1/B[19] ), .A2(\intadd_1/A[19] ), .ZN(
        \intadd_1/n64 ) );
  AOI21_X1 U4528 ( .B1(n5325), .B2(n4247), .A(n7211), .ZN(\intadd_1/B[19] ) );
  AOI21_X1 U4529 ( .B1(\intadd_1/n140 ), .B2(\intadd_1/n91 ), .A(
        \intadd_1/n92 ), .ZN(\intadd_1/n90 ) );
  OAI21_X1 U4530 ( .B1(\intadd_1/n119 ), .B2(\intadd_1/n93 ), .A(
        \intadd_1/n94 ), .ZN(\intadd_1/n92 ) );
  OAI21_X1 U4531 ( .B1(\intadd_1/n138 ), .B2(\intadd_1/n134 ), .A(
        \intadd_1/n135 ), .ZN(n4720) );
  OAI21_X1 U4532 ( .B1(\intadd_1/n161 ), .B2(\intadd_1/n141 ), .A(
        \intadd_1/n142 ), .ZN(\intadd_1/n140 ) );
  AOI21_X1 U4533 ( .B1(n4029), .B2(\intadd_1/n162 ), .A(\intadd_1/n163 ), .ZN(
        \intadd_1/n161 ) );
  NOR2_X1 U4534 ( .A1(n5272), .A2(n7247), .ZN(\intadd_1/A[1] ) );
  NOR2_X1 U4535 ( .A1(\intadd_1/A[2] ), .A2(\intadd_1/B[2] ), .ZN(
        \intadd_1/n164 ) );
  NOR2_X1 U4536 ( .A1(n5322), .A2(n7245), .ZN(\intadd_1/B[2] ) );
  NOR2_X1 U4537 ( .A1(\intadd_1/n148 ), .A2(\intadd_1/n145 ), .ZN(
        \intadd_1/n143 ) );
  NOR2_X1 U4538 ( .A1(\intadd_1/A[5] ), .A2(\intadd_1/B[5] ), .ZN(
        \intadd_1/n148 ) );
  AOI21_X1 U4539 ( .B1(n5325), .B2(n4254), .A(n7239), .ZN(\intadd_1/B[5] ) );
  XNOR2_X1 U4540 ( .A(n5865), .B(sub_add_exe), .ZN(\intadd_1/A[5] ) );
  AOI21_X1 U4541 ( .B1(n3903), .B2(n4340), .A(n5259), .ZN(n5865) );
  AOI21_X1 U4542 ( .B1(n5118), .B2(n4253), .A(n7237), .ZN(\intadd_1/B[6] ) );
  NOR2_X1 U4543 ( .A1(\intadd_1/n153 ), .A2(\intadd_1/n158 ), .ZN(
        \intadd_1/n151 ) );
  NOR2_X1 U4544 ( .A1(\intadd_1/A[3] ), .A2(\intadd_1/B[3] ), .ZN(
        \intadd_1/n158 ) );
  NOR2_X1 U4545 ( .A1(n5320), .A2(n7243), .ZN(\intadd_1/B[3] ) );
  NOR2_X1 U4546 ( .A1(n4668), .A2(\intadd_1/B[4] ), .ZN(\intadd_1/n153 ) );
  OAI211_X1 U4547 ( .C1(n4671), .C2(n4734), .A(n4670), .B(n4669), .ZN(n4668)
         );
  AND2_X1 U4548 ( .A1(n3903), .A2(n4330), .ZN(n4734) );
  NOR2_X1 U4549 ( .A1(\intadd_1/n118 ), .A2(\intadd_1/n93 ), .ZN(
        \intadd_1/n91 ) );
  NAND2_X1 U4550 ( .A1(\intadd_1/n95 ), .A2(\intadd_1/n107 ), .ZN(
        \intadd_1/n93 ) );
  NOR2_X1 U4551 ( .A1(\intadd_1/n102 ), .A2(\intadd_1/n97 ), .ZN(
        \intadd_1/n95 ) );
  NOR2_X1 U4552 ( .A1(n5302), .A2(n7221), .ZN(\intadd_1/B[14] ) );
  XNOR2_X1 U4553 ( .A(n5116), .B(sub_add_exe), .ZN(\intadd_1/A[14] ) );
  NOR2_X1 U4554 ( .A1(\intadd_1/A[13] ), .A2(\intadd_1/B[13] ), .ZN(
        \intadd_1/n102 ) );
  AOI21_X1 U4555 ( .B1(n5118), .B2(n4250), .A(n7223), .ZN(\intadd_1/B[13] ) );
  XNOR2_X1 U4556 ( .A(n5012), .B(sub_add_exe), .ZN(\intadd_1/A[13] ) );
  AOI21_X1 U4557 ( .B1(n5119), .B2(n4306), .A(n5250), .ZN(n5012) );
  NOR2_X1 U4558 ( .A1(\intadd_1/n114 ), .A2(\intadd_1/n109 ), .ZN(
        \intadd_1/n107 ) );
  AOI21_X1 U4559 ( .B1(n5325), .B2(n4251), .A(n7225), .ZN(\intadd_1/B[12] ) );
  XNOR2_X1 U4560 ( .A(n4938), .B(n4225), .ZN(\intadd_1/A[12] ) );
  NOR2_X1 U4561 ( .A1(\intadd_1/A[11] ), .A2(\intadd_1/B[11] ), .ZN(
        \intadd_1/n114 ) );
  AOI21_X1 U4562 ( .B1(n5325), .B2(n4252), .A(n7227), .ZN(\intadd_1/B[11] ) );
  XNOR2_X1 U4563 ( .A(n5005), .B(sub_add_exe), .ZN(\intadd_1/A[11] ) );
  AOI21_X1 U4564 ( .B1(n5122), .B2(n4305), .A(n5252), .ZN(n5005) );
  NAND2_X1 U4565 ( .A1(\intadd_1/n120 ), .A2(\intadd_1/n132 ), .ZN(
        \intadd_1/n118 ) );
  NOR2_X1 U4566 ( .A1(\intadd_1/n137 ), .A2(\intadd_1/n134 ), .ZN(
        \intadd_1/n132 ) );
  NOR2_X1 U4567 ( .A1(n5313), .A2(n7233), .ZN(\intadd_1/B[8] ) );
  OAI21_X1 U4568 ( .B1(n4705), .B2(\dp/b_adder_id_exe_int[9] ), .A(n5256), 
        .ZN(n5144) );
  NOR2_X1 U4569 ( .A1(\intadd_1/B[7] ), .A2(\intadd_1/A[7] ), .ZN(
        \intadd_1/n137 ) );
  XNOR2_X1 U4570 ( .A(n5894), .B(n4225), .ZN(\intadd_1/A[7] ) );
  NAND2_X1 U4571 ( .A1(n5258), .A2(n5257), .ZN(n5894) );
  NOR2_X1 U4572 ( .A1(n7235), .A2(n5315), .ZN(\intadd_1/B[7] ) );
  NOR2_X1 U4573 ( .A1(n4038), .A2(\intadd_1/B[10] ), .ZN(n4706) );
  NOR2_X1 U4574 ( .A1(n7229), .A2(n5309), .ZN(\intadd_1/B[10] ) );
  NOR2_X1 U4575 ( .A1(\intadd_1/A[9] ), .A2(\intadd_1/B[9] ), .ZN(
        \intadd_1/n127 ) );
  NOR2_X1 U4576 ( .A1(n7231), .A2(n5311), .ZN(\intadd_1/B[9] ) );
  OR2_X1 U4577 ( .A1(\intadd_1/A[25] ), .A2(\intadd_1/B[25] ), .ZN(n4229) );
  AOI21_X1 U4578 ( .B1(n5118), .B2(n4241), .A(n7199), .ZN(\intadd_1/B[25] ) );
  XNOR2_X1 U4579 ( .A(n6082), .B(sub_add_exe), .ZN(\intadd_1/A[25] ) );
  AOI21_X1 U4580 ( .B1(n5170), .B2(n4291), .A(n5240), .ZN(n6082) );
  AND2_X1 U4581 ( .A1(\intadd_1/n37 ), .A2(n4776), .ZN(n4352) );
  OR2_X1 U4582 ( .A1(\intadd_1/A[26] ), .A2(\intadd_1/B[26] ), .ZN(n4776) );
  NOR2_X1 U4583 ( .A1(n5285), .A2(n7197), .ZN(\intadd_1/B[26] ) );
  XNOR2_X1 U4584 ( .A(n6096), .B(n4225), .ZN(\intadd_1/A[26] ) );
  AOI21_X1 U4585 ( .B1(n5118), .B2(n4242), .A(n7201), .ZN(\intadd_1/B[24] ) );
  INV_X1 U4586 ( .A(n5081), .ZN(n4797) );
  INV_X1 U4587 ( .A(n7253), .ZN(n5325) );
  AND2_X1 U4588 ( .A1(n5264), .A2(\ctrl_u/curr_mem[3] ), .ZN(n5266) );
  XNOR2_X1 U4589 ( .A(rs_exe[0]), .B(rd_exemem[0]), .ZN(n5264) );
  XNOR2_X1 U4590 ( .A(n6065), .B(n4225), .ZN(\intadd_1/A[24] ) );
  AND2_X2 U4591 ( .A1(n4022), .A2(n5061), .ZN(n4726) );
  NOR2_X1 U4592 ( .A1(n5141), .A2(n5139), .ZN(n5135) );
  NAND2_X1 U4593 ( .A1(n5342), .A2(n4300), .ZN(n4738) );
  NAND2_X1 U4594 ( .A1(n4840), .A2(n4728), .ZN(n5342) );
  AND2_X1 U4595 ( .A1(n4959), .A2(n4842), .ZN(n4840) );
  NAND4_X1 U4596 ( .A1(n4742), .A2(n4022), .A3(n4739), .A4(n4741), .ZN(n5768)
         );
  NAND2_X1 U4597 ( .A1(n5062), .A2(n4740), .ZN(n4739) );
  NOR2_X1 U4598 ( .A1(n4743), .A2(n4744), .ZN(n4742) );
  AND4_X2 U4599 ( .A1(n5098), .A2(n4232), .A3(n3924), .A4(n4839), .ZN(n5141)
         );
  AND2_X1 U4600 ( .A1(n5061), .A2(n4300), .ZN(n4839) );
  NAND2_X1 U4601 ( .A1(n4318), .A2(n7273), .ZN(n4799) );
  NAND2_X1 U4602 ( .A1(n4015), .A2(\ctrl_u/curr_ms ), .ZN(n4703) );
  XNOR2_X1 U4603 ( .A(rt_exe[1]), .B(rd_exemem[1]), .ZN(n4960) );
  XNOR2_X1 U4604 ( .A(rt_exe[0]), .B(rd_exemem[0]), .ZN(n5239) );
  XNOR2_X1 U4605 ( .A(rt_exe[3]), .B(rd_exemem[3]), .ZN(n4841) );
  OR2_X1 U4606 ( .A1(n5173), .A2(n4109), .ZN(n5276) );
  NOR2_X1 U4607 ( .A1(n5174), .A2(n493), .ZN(n5277) );
  NAND2_X1 U4608 ( .A1(n5657), .A2(n5670), .ZN(n5668) );
  AND2_X1 U4609 ( .A1(n4711), .A2(n4710), .ZN(n4836) );
  AND2_X1 U4610 ( .A1(n4841), .A2(n4842), .ZN(n4736) );
  OR2_X1 U4611 ( .A1(n6315), .A2(n6510), .ZN(n6534) );
  NOR2_X1 U4612 ( .A1(op_b_fw_sel_exe[1]), .A2(n7444), .ZN(n7445) );
  INV_X1 U4613 ( .A(n5165), .ZN(n5155) );
  NOR2_X1 U4614 ( .A1(n5026), .A2(n5229), .ZN(n5025) );
  OAI21_X1 U4615 ( .B1(n7312), .B2(n5413), .A(n5389), .ZN(n6333) );
  NOR2_X1 U4616 ( .A1(n5668), .A2(n3924), .ZN(n5389) );
  OR2_X1 U4617 ( .A1(n5655), .A2(\ctrl_u/N1805 ), .ZN(n5657) );
  INV_X1 U4618 ( .A(n7445), .ZN(n7446) );
  AND2_X1 U4619 ( .A1(n6480), .A2(n6477), .ZN(n6486) );
  INV_X1 U4620 ( .A(wp_data[30]), .ZN(n5274) );
  OR2_X1 U4621 ( .A1(n5173), .A2(n4068), .ZN(n5280) );
  NOR2_X1 U4622 ( .A1(\ctrl_u/curr_exe_39 ), .A2(\ctrl_u/curr_exe_40 ), .ZN(
        n5671) );
  OR2_X1 U4623 ( .A1(\dp/b10_1_mult_id_exe_int[1] ), .A2(n593), .ZN(n5681) );
  INV_X1 U4624 ( .A(n5148), .ZN(n5149) );
  NOR2_X1 U4625 ( .A1(pc_en), .A2(n5229), .ZN(n7108) );
  NOR2_X1 U4626 ( .A1(en_b_exe), .A2(n7442), .ZN(n7492) );
  NAND2_X1 U4627 ( .A1(n4762), .A2(\ctrl_u/curr_mul_in_prog ), .ZN(n5234) );
  INV_X1 U4628 ( .A(n6334), .ZN(n4921) );
  BUF_X2 U4629 ( .A(n5156), .Z(n5186) );
  BUF_X2 U4630 ( .A(n6298), .Z(n5189) );
  NAND2_X1 U4631 ( .A1(\ctrl_u/mem_stall ), .A2(\ctrl_u/curr_ak_exe ), .ZN(
        n5337) );
  NOR2_X1 U4632 ( .A1(n7089), .A2(alu_comp_sel[0]), .ZN(n5754) );
  NOR2_X1 U4633 ( .A1(n7146), .A2(b_selector_id), .ZN(n6980) );
  OR2_X1 U4634 ( .A1(n5618), .A2(n7312), .ZN(n4237) );
  XNOR2_X1 U4635 ( .A(\dp/npc_id_exe_int[3] ), .B(\dp/npc_id_exe_int[2] ), 
        .ZN(btb_cache_rw_address[1]) );
  NAND2_X1 U4636 ( .A1(n6175), .A2(n6174), .ZN(btb_cache_rw_address[2]) );
  INV_X1 U4637 ( .A(n7370), .ZN(n6174) );
  OAI21_X1 U4638 ( .B1(\dp/npc_id_exe_int[2] ), .B2(\dp/npc_id_exe_int[3] ), 
        .A(\dp/npc_id_exe_int[4] ), .ZN(n6175) );
  NOR3_X1 U4639 ( .A1(\dp/npc_id_exe_int[3] ), .A2(\dp/npc_id_exe_int[4] ), 
        .A3(\dp/npc_id_exe_int[2] ), .ZN(n7370) );
  OAI21_X1 U4640 ( .B1(n5810), .B2(n7526), .A(n5774), .ZN(ram_data_in[4]) );
  NAND2_X1 U4641 ( .A1(n5191), .A2(n4610), .ZN(n5774) );
  OAI21_X1 U4642 ( .B1(n5810), .B2(n7522), .A(n5772), .ZN(ram_data_in[2]) );
  NAND2_X1 U4643 ( .A1(n5810), .A2(n4608), .ZN(n5772) );
  OAI21_X1 U4644 ( .B1(n5190), .B2(n7528), .A(n5776), .ZN(ram_data_in[6]) );
  NAND2_X1 U4645 ( .A1(n5810), .A2(n4612), .ZN(n5776) );
  OAI21_X1 U4646 ( .B1(n5191), .B2(n7502), .A(n5781), .ZN(ram_data_in[11]) );
  NAND2_X1 U4647 ( .A1(n5191), .A2(n4617), .ZN(n5781) );
  OAI21_X1 U4648 ( .B1(n5191), .B2(n7503), .A(n5782), .ZN(ram_data_in[12]) );
  NAND2_X1 U4649 ( .A1(n5191), .A2(n4618), .ZN(n5782) );
  OAI21_X1 U4650 ( .B1(n5810), .B2(n7525), .A(n5773), .ZN(ram_data_in[3]) );
  NAND2_X1 U4651 ( .A1(n5810), .A2(n4609), .ZN(n5773) );
  OAI21_X1 U4652 ( .B1(n5190), .B2(n7531), .A(n5779), .ZN(ram_data_in[9]) );
  NAND2_X1 U4653 ( .A1(n5810), .A2(n4615), .ZN(n5779) );
  OAI21_X1 U4654 ( .B1(n5190), .B2(n7523), .A(n5800), .ZN(ram_data_in[30]) );
  NAND2_X1 U4655 ( .A1(n5191), .A2(n4636), .ZN(n5800) );
  OAI21_X1 U4656 ( .B1(n5190), .B2(n7530), .A(n5778), .ZN(ram_data_in[8]) );
  NAND2_X1 U4657 ( .A1(n5810), .A2(n4614), .ZN(n5778) );
  OAI21_X1 U4658 ( .B1(n5190), .B2(n7529), .A(n5777), .ZN(ram_data_in[7]) );
  NAND2_X1 U4659 ( .A1(n5810), .A2(n4613), .ZN(n5777) );
  OAI21_X1 U4660 ( .B1(n5190), .B2(n7507), .A(n5786), .ZN(ram_data_in[16]) );
  NAND2_X1 U4661 ( .A1(n5191), .A2(n4622), .ZN(n5786) );
  OAI21_X1 U4662 ( .B1(n5191), .B2(n7510), .A(n5789), .ZN(ram_data_in[19]) );
  NAND2_X1 U4663 ( .A1(n5191), .A2(n4625), .ZN(n5789) );
  OAI21_X1 U4664 ( .B1(n5810), .B2(n7527), .A(n5775), .ZN(ram_data_in[5]) );
  NAND2_X1 U4665 ( .A1(n5810), .A2(n4611), .ZN(n5775) );
  OAI21_X1 U4666 ( .B1(n5191), .B2(n7524), .A(n5801), .ZN(ram_data_in[31]) );
  NAND2_X1 U4667 ( .A1(n5191), .A2(n4637), .ZN(n5801) );
  OAI21_X1 U4668 ( .B1(n5191), .B2(n7521), .A(n5799), .ZN(ram_data_in[29]) );
  NAND2_X1 U4669 ( .A1(n5810), .A2(n4635), .ZN(n5799) );
  OAI21_X1 U4670 ( .B1(n5191), .B2(n7520), .A(n5798), .ZN(ram_data_in[28]) );
  NAND2_X1 U4671 ( .A1(n5810), .A2(n4634), .ZN(n5798) );
  OAI21_X1 U4672 ( .B1(n5191), .B2(n7519), .A(n5797), .ZN(ram_data_in[27]) );
  NAND2_X1 U4673 ( .A1(n5191), .A2(n4633), .ZN(n5797) );
  OAI21_X1 U4674 ( .B1(n5191), .B2(n7518), .A(n5796), .ZN(ram_data_in[26]) );
  NAND2_X1 U4675 ( .A1(n5191), .A2(n4632), .ZN(n5796) );
  OAI21_X1 U4676 ( .B1(n5810), .B2(n7511), .A(n5771), .ZN(ram_data_in[1]) );
  NAND2_X1 U4677 ( .A1(n5191), .A2(n4607), .ZN(n5771) );
  OAI21_X1 U4678 ( .B1(n5810), .B2(n7500), .A(n5770), .ZN(ram_data_in[0]) );
  NAND2_X1 U4679 ( .A1(n5810), .A2(n4606), .ZN(n5770) );
  OAI21_X1 U4680 ( .B1(n5191), .B2(n7501), .A(n5780), .ZN(ram_data_in[10]) );
  NAND2_X1 U4681 ( .A1(n5191), .A2(n4616), .ZN(n5780) );
  OAI21_X1 U4682 ( .B1(n5810), .B2(n7517), .A(n5795), .ZN(ram_data_in[25]) );
  NAND2_X1 U4683 ( .A1(n5191), .A2(n4631), .ZN(n5795) );
  OAI21_X1 U4684 ( .B1(n5810), .B2(n7516), .A(n5794), .ZN(ram_data_in[24]) );
  NAND2_X1 U4685 ( .A1(n5191), .A2(n4630), .ZN(n5794) );
  OAI21_X1 U4686 ( .B1(n5810), .B2(n7515), .A(n5793), .ZN(ram_data_in[23]) );
  NAND2_X1 U4687 ( .A1(n5191), .A2(n4629), .ZN(n5793) );
  OAI21_X1 U4688 ( .B1(n5191), .B2(n7514), .A(n5792), .ZN(ram_data_in[22]) );
  NAND2_X1 U4689 ( .A1(n5191), .A2(n4628), .ZN(n5792) );
  OAI21_X1 U4690 ( .B1(n5191), .B2(n7513), .A(n5791), .ZN(ram_data_in[21]) );
  NAND2_X1 U4691 ( .A1(n5191), .A2(n4627), .ZN(n5791) );
  OAI21_X1 U4692 ( .B1(n5191), .B2(n7512), .A(n5790), .ZN(ram_data_in[20]) );
  NAND2_X1 U4693 ( .A1(n5191), .A2(n4626), .ZN(n5790) );
  OAI21_X1 U4694 ( .B1(n5810), .B2(n7506), .A(n5785), .ZN(ram_data_in[15]) );
  NAND2_X1 U4695 ( .A1(n5191), .A2(n4621), .ZN(n5785) );
  OAI21_X1 U4696 ( .B1(n5191), .B2(n7509), .A(n5788), .ZN(ram_data_in[18]) );
  NAND2_X1 U4697 ( .A1(n5810), .A2(n4624), .ZN(n5788) );
  OAI21_X1 U4698 ( .B1(n5191), .B2(n7508), .A(n5787), .ZN(ram_data_in[17]) );
  NAND2_X1 U4699 ( .A1(n5810), .A2(n4623), .ZN(n5787) );
  OAI21_X1 U4700 ( .B1(n5191), .B2(n7505), .A(n5784), .ZN(ram_data_in[14]) );
  NAND2_X1 U4701 ( .A1(n5810), .A2(n4620), .ZN(n5784) );
  OAI21_X1 U4702 ( .B1(n5190), .B2(n7504), .A(n5783), .ZN(ram_data_in[13]) );
  NAND2_X1 U4703 ( .A1(n5191), .A2(n4619), .ZN(n5783) );
  OR2_X1 U4704 ( .A1(n5753), .A2(n5229), .ZN(\ctrl_u/n560 ) );
  INV_X1 U4705 ( .A(n5807), .ZN(ram_address[5]) );
  AOI222_X1 U4706 ( .A1(n4643), .A2(n5191), .B1(ram_rw), .B2(
        cpu_cache_address[5]), .C1(n5809), .C2(evicted_cache_address[5]), .ZN(
        n5807) );
  INV_X1 U4707 ( .A(n5811), .ZN(ram_address[7]) );
  AOI222_X1 U4708 ( .A1(n4645), .A2(n5191), .B1(ram_rw), .B2(
        cpu_cache_address[7]), .C1(n5809), .C2(evicted_cache_address[7]), .ZN(
        n5811) );
  INV_X1 U4709 ( .A(n5805), .ZN(ram_address[3]) );
  AOI222_X1 U4710 ( .A1(n4641), .A2(n5190), .B1(ram_rw), .B2(
        cpu_cache_address[3]), .C1(n5809), .C2(evicted_cache_address[3]), .ZN(
        n5805) );
  INV_X1 U4711 ( .A(n5808), .ZN(ram_address[6]) );
  AOI222_X1 U4712 ( .A1(n4644), .A2(n5191), .B1(ram_rw), .B2(
        cpu_cache_address[6]), .C1(n5809), .C2(evicted_cache_address[6]), .ZN(
        n5808) );
  INV_X1 U4713 ( .A(n5803), .ZN(ram_address[1]) );
  AOI222_X1 U4714 ( .A1(n4639), .A2(n5190), .B1(ram_rw), .B2(
        cpu_cache_address[1]), .C1(n5809), .C2(evicted_cache_address[1]), .ZN(
        n5803) );
  INV_X1 U4715 ( .A(n5802), .ZN(ram_address[0]) );
  AOI222_X1 U4716 ( .A1(n4638), .A2(n5190), .B1(ram_rw), .B2(
        cpu_cache_address[0]), .C1(n5809), .C2(evicted_cache_address[0]), .ZN(
        n5802) );
  INV_X1 U4717 ( .A(n5804), .ZN(ram_address[2]) );
  AOI222_X1 U4718 ( .A1(n4640), .A2(n5190), .B1(ram_rw), .B2(
        cpu_cache_address[2]), .C1(n5809), .C2(evicted_cache_address[2]), .ZN(
        n5804) );
  INV_X1 U4719 ( .A(n5806), .ZN(ram_address[4]) );
  AOI222_X1 U4720 ( .A1(n4642), .A2(n5191), .B1(ram_rw), .B2(
        cpu_cache_address[4]), .C1(n5809), .C2(evicted_cache_address[4]), .ZN(
        n5806) );
  NOR2_X1 U4721 ( .A1(n5190), .A2(n5809), .ZN(ram_rw) );
  NAND2_X1 U4722 ( .A1(n5665), .A2(n5662), .ZN(\ctrl_u/next_mem[3] ) );
  NAND2_X1 U4723 ( .A1(n5665), .A2(n5663), .ZN(\ctrl_u/next_mem[4] ) );
  NAND2_X1 U4724 ( .A1(n5665), .A2(n5661), .ZN(\ctrl_u/next_mem[2] ) );
  NAND2_X1 U4725 ( .A1(n5665), .A2(n5664), .ZN(\ctrl_u/next_mem[6] ) );
  NOR2_X1 U4726 ( .A1(n5669), .A2(n5660), .ZN(n5665) );
  INV_X1 U4727 ( .A(rst_exe_mem_regs), .ZN(n5660) );
  NAND2_X1 U4728 ( .A1(ram_update), .A2(rst_mem_wb_regs), .ZN(n5678) );
  OAI22_X1 U4729 ( .A1(n5666), .A2(n4180), .B1(n5670), .B2(n4479), .ZN(
        \ctrl_u/next_mem[7] ) );
  OAI22_X1 U4730 ( .A1(n5666), .A2(n4181), .B1(n5670), .B2(n4470), .ZN(
        \ctrl_u/next_mem[8] ) );
  OAI22_X1 U4731 ( .A1(n5666), .A2(n4450), .B1(n5670), .B2(n4166), .ZN(
        \ctrl_u/next_mem[10] ) );
  INV_X1 U4732 ( .A(n5667), .ZN(n5666) );
  AOI21_X1 U4733 ( .B1(n5656), .B2(n5672), .A(n5668), .ZN(n5667) );
  INV_X1 U4734 ( .A(n5659), .ZN(n5656) );
  OAI21_X1 U4735 ( .B1(n7392), .B2(n4525), .A(n7386), .ZN(n3136) );
  OAI21_X1 U4736 ( .B1(n7392), .B2(n4524), .A(n7385), .ZN(n3137) );
  OAI21_X1 U4737 ( .B1(n7392), .B2(n4526), .A(n7387), .ZN(n3135) );
  OAI21_X1 U4738 ( .B1(n7392), .B2(n4523), .A(n7384), .ZN(n3138) );
  OAI21_X1 U4739 ( .B1(n7392), .B2(n4527), .A(n7388), .ZN(n3134) );
  OAI21_X1 U4740 ( .B1(n7392), .B2(n4529), .A(n7390), .ZN(n3132) );
  OAI21_X1 U4741 ( .B1(n7392), .B2(n4528), .A(n7389), .ZN(n3133) );
  OAI211_X1 U4742 ( .C1(n7392), .C2(n4538), .A(n7393), .B(n7391), .ZN(n3131)
         );
  OAI222_X1 U4743 ( .A1(n4096), .A2(n7497), .B1(n7498), .B2(n4436), .C1(n4149), 
        .C2(n7499), .ZN(n2558) );
  OAI222_X1 U4744 ( .A1(n4506), .A2(n7498), .B1(n4081), .B2(n7497), .C1(n4150), 
        .C2(n7499), .ZN(n2574) );
  OAI222_X1 U4745 ( .A1(n4512), .A2(n7498), .B1(n4082), .B2(n7497), .C1(n4156), 
        .C2(n7499), .ZN(n2580) );
  OAI222_X1 U4746 ( .A1(n4514), .A2(n7498), .B1(n6453), .B2(n7497), .C1(n4158), 
        .C2(n7499), .ZN(n2582) );
  OAI222_X1 U4747 ( .A1(n4109), .A2(n7497), .B1(n7496), .B2(n7498), .C1(n4401), 
        .C2(n7499), .ZN(n2559) );
  OAI222_X1 U4748 ( .A1(n4080), .A2(n7497), .B1(n7498), .B2(n4438), .C1(n4162), 
        .C2(n7499), .ZN(n2586) );
  OAI222_X1 U4749 ( .A1(n4071), .A2(n7497), .B1(n7498), .B2(n4437), .C1(n4161), 
        .C2(n7499), .ZN(n2585) );
  OAI222_X1 U4750 ( .A1(n4377), .A2(n7497), .B1(n7498), .B2(n4440), .C1(n4164), 
        .C2(n7499), .ZN(n2589) );
  OAI222_X1 U4751 ( .A1(n4072), .A2(n7497), .B1(n7498), .B2(n4439), .C1(n4163), 
        .C2(n7499), .ZN(n2588) );
  OAI222_X1 U4752 ( .A1(n4087), .A2(n7497), .B1(n7498), .B2(n4441), .C1(n4165), 
        .C2(n7499), .ZN(n2587) );
  OAI222_X1 U4753 ( .A1(n4516), .A2(n7498), .B1(n6459), .B2(n7497), .C1(n4160), 
        .C2(n7499), .ZN(n2584) );
  OAI222_X1 U4754 ( .A1(n4515), .A2(n7498), .B1(n6456), .B2(n7497), .C1(n4159), 
        .C2(n7499), .ZN(n2583) );
  AOI22_X1 U4755 ( .A1(n3958), .A2(wp_data[17]), .B1(dcache_data_out[17]), 
        .B2(n3959), .ZN(n7465) );
  AOI22_X1 U4756 ( .A1(n3958), .A2(wp_data[21]), .B1(dcache_data_out[21]), 
        .B2(n7492), .ZN(n7473) );
  AOI22_X1 U4757 ( .A1(n3958), .A2(wp_data[18]), .B1(dcache_data_out[18]), 
        .B2(n3959), .ZN(n7467) );
  AOI22_X1 U4758 ( .A1(n3958), .A2(wp_data[23]), .B1(dcache_data_out[23]), 
        .B2(n7492), .ZN(n7477) );
  AOI22_X1 U4759 ( .A1(n3958), .A2(wp_data[22]), .B1(dcache_data_out[22]), 
        .B2(n3959), .ZN(n7475) );
  AOI22_X1 U4760 ( .A1(n3958), .A2(wp_data[20]), .B1(dcache_data_out[20]), 
        .B2(n3959), .ZN(n7471) );
  AOI22_X1 U4761 ( .A1(n3958), .A2(wp_data[19]), .B1(dcache_data_out[19]), 
        .B2(n3959), .ZN(n7469) );
  AOI22_X1 U4762 ( .A1(n3958), .A2(wp_data[28]), .B1(n3959), .B2(
        dcache_data_out[28]), .ZN(n7487) );
  AOI22_X1 U4763 ( .A1(n3958), .A2(wp_data[24]), .B1(n3959), .B2(
        dcache_data_out[24]), .ZN(n7479) );
  AOI22_X1 U4764 ( .A1(n3958), .A2(wp_data[29]), .B1(n3959), .B2(
        dcache_data_out[29]), .ZN(n7489) );
  AOI22_X1 U4765 ( .A1(n3958), .A2(wp_data[27]), .B1(n3959), .B2(
        dcache_data_out[27]), .ZN(n7485) );
  AOI22_X1 U4766 ( .A1(n3958), .A2(wp_data[25]), .B1(n3959), .B2(
        dcache_data_out[25]), .ZN(n7481) );
  AOI22_X1 U4767 ( .A1(n3958), .A2(wp_data[26]), .B1(n7492), .B2(
        dcache_data_out[26]), .ZN(n7483) );
  OAI211_X1 U4768 ( .C1(n7495), .C2(n4088), .A(n7459), .B(n6441), .ZN(n2609)
         );
  AOI22_X1 U4769 ( .A1(n3958), .A2(wp_data[12]), .B1(dcache_data_out[12]), 
        .B2(n3959), .ZN(n6441) );
  OAI211_X1 U4770 ( .C1(n7495), .C2(n4087), .A(n7449), .B(n7099), .ZN(n2619)
         );
  AOI22_X1 U4771 ( .A1(n3958), .A2(wp_data[2]), .B1(dcache_data_out[2]), .B2(
        n3959), .ZN(n7099) );
  OAI211_X1 U4772 ( .C1(n7495), .C2(n4066), .A(n7461), .B(n6435), .ZN(n2607)
         );
  AOI22_X1 U4773 ( .A1(n3958), .A2(wp_data[14]), .B1(dcache_data_out[14]), 
        .B2(n3959), .ZN(n6435) );
  OAI211_X1 U4774 ( .C1(n7495), .C2(n4377), .A(n7447), .B(n6185), .ZN(n2621)
         );
  AOI22_X1 U4775 ( .A1(n3958), .A2(wp_data[0]), .B1(dcache_data_out[0]), .B2(
        n3959), .ZN(n6185) );
  OAI211_X1 U4776 ( .C1(n7495), .C2(n4081), .A(n7462), .B(n6433), .ZN(n2606)
         );
  AOI22_X1 U4777 ( .A1(n3958), .A2(wp_data[15]), .B1(dcache_data_out[15]), 
        .B2(n3959), .ZN(n6433) );
  OAI211_X1 U4778 ( .C1(n7495), .C2(n4082), .A(n7456), .B(n6448), .ZN(n2612)
         );
  AOI22_X1 U4779 ( .A1(n3958), .A2(wp_data[9]), .B1(dcache_data_out[9]), .B2(
        n3959), .ZN(n6448) );
  OAI211_X1 U4780 ( .C1(n7495), .C2(n4073), .A(n7458), .B(n6444), .ZN(n2610)
         );
  AOI22_X1 U4781 ( .A1(n3958), .A2(wp_data[11]), .B1(dcache_data_out[11]), 
        .B2(n3959), .ZN(n6444) );
  OAI211_X1 U4782 ( .C1(n7495), .C2(n4079), .A(n7460), .B(n6438), .ZN(n2608)
         );
  AOI22_X1 U4783 ( .A1(n3958), .A2(wp_data[13]), .B1(dcache_data_out[13]), 
        .B2(n3959), .ZN(n6438) );
  OAI211_X1 U4784 ( .C1(n7495), .C2(n4074), .A(n7457), .B(n6446), .ZN(n2611)
         );
  AOI22_X1 U4785 ( .A1(n3958), .A2(wp_data[10]), .B1(dcache_data_out[10]), 
        .B2(n3959), .ZN(n6446) );
  OAI211_X1 U4786 ( .C1(n7495), .C2(n4071), .A(n7451), .B(n6461), .ZN(n2617)
         );
  AOI22_X1 U4787 ( .A1(n3958), .A2(wp_data[4]), .B1(dcache_data_out[4]), .B2(
        n3959), .ZN(n6461) );
  OAI211_X1 U4788 ( .C1(n7495), .C2(n4109), .A(n7490), .B(n6411), .ZN(n2591)
         );
  AOI22_X1 U4789 ( .A1(n3958), .A2(wp_data[30]), .B1(n7492), .B2(
        dcache_data_out[30]), .ZN(n6411) );
  OAI211_X1 U4790 ( .C1(n7495), .C2(n4089), .A(n7463), .B(n6432), .ZN(n2605)
         );
  AOI22_X1 U4791 ( .A1(n3958), .A2(wp_data[16]), .B1(dcache_data_out[16]), 
        .B2(n3959), .ZN(n6432) );
  OAI211_X1 U4792 ( .C1(n7495), .C2(n6453), .A(n7454), .B(n6452), .ZN(n2614)
         );
  AOI22_X1 U4793 ( .A1(n3958), .A2(wp_data[7]), .B1(dcache_data_out[7]), .B2(
        n3959), .ZN(n6452) );
  OAI211_X1 U4794 ( .C1(n7495), .C2(n4080), .A(n7450), .B(n6463), .ZN(n2618)
         );
  AOI22_X1 U4795 ( .A1(n3958), .A2(wp_data[3]), .B1(dcache_data_out[3]), .B2(
        n3959), .ZN(n6463) );
  OAI211_X1 U4796 ( .C1(n7495), .C2(n4072), .A(n7448), .B(n6465), .ZN(n2620)
         );
  AOI22_X1 U4797 ( .A1(n3958), .A2(wp_data[1]), .B1(dcache_data_out[1]), .B2(
        n3959), .ZN(n6465) );
  OAI211_X1 U4798 ( .C1(n7495), .C2(n4096), .A(n7494), .B(n6335), .ZN(n2590)
         );
  AOI22_X1 U4799 ( .A1(n3958), .A2(wp_data[31]), .B1(dcache_data_out[31]), 
        .B2(n3959), .ZN(n6335) );
  OAI211_X1 U4800 ( .C1(n7495), .C2(n4063), .A(n7455), .B(n6450), .ZN(n2613)
         );
  AOI22_X1 U4801 ( .A1(n3958), .A2(wp_data[8]), .B1(dcache_data_out[8]), .B2(
        n3959), .ZN(n6450) );
  OAI211_X1 U4802 ( .C1(n7495), .C2(n6456), .A(n7453), .B(n6455), .ZN(n2615)
         );
  AOI22_X1 U4803 ( .A1(n3958), .A2(wp_data[6]), .B1(dcache_data_out[6]), .B2(
        n3959), .ZN(n6455) );
  OAI211_X1 U4804 ( .C1(n7495), .C2(n6459), .A(n7452), .B(n6458), .ZN(n2616)
         );
  AOI22_X1 U4805 ( .A1(n3958), .A2(wp_data[5]), .B1(dcache_data_out[5]), .B2(
        n3959), .ZN(n6458) );
  OR2_X1 U4806 ( .A1(n5657), .A2(n7340), .ZN(rst_exe_mem_regs) );
  INV_X1 U4807 ( .A(n5342), .ZN(n5767) );
  OAI222_X1 U4808 ( .A1(n4513), .A2(n7498), .B1(n4063), .B2(n7497), .C1(n4157), 
        .C2(n7499), .ZN(n2581) );
  OAI222_X1 U4809 ( .A1(n4507), .A2(n7498), .B1(n4066), .B2(n7497), .C1(n4151), 
        .C2(n7499), .ZN(n2575) );
  OAI222_X1 U4810 ( .A1(n4511), .A2(n7498), .B1(n4074), .B2(n7497), .C1(n4155), 
        .C2(n7499), .ZN(n2579) );
  OAI222_X1 U4811 ( .A1(n4508), .A2(n7498), .B1(n4079), .B2(n7497), .C1(n4152), 
        .C2(n7499), .ZN(n2576) );
  OAI222_X1 U4812 ( .A1(n4510), .A2(n7498), .B1(n4073), .B2(n7497), .C1(n4154), 
        .C2(n7499), .ZN(n2578) );
  OAI222_X1 U4813 ( .A1(n4509), .A2(n7498), .B1(n4088), .B2(n7497), .C1(n4153), 
        .C2(n7499), .ZN(n2577) );
  OAI22_X1 U4814 ( .A1(n6447), .A2(n7440), .B1(n4074), .B2(n3938), .ZN(n2643)
         );
  OAI21_X1 U4815 ( .B1(n6173), .B2(btb_cache_data_out_rw[30]), .A(n6170), .ZN(
        btb_cache_data_in[30]) );
  OAI211_X1 U4816 ( .C1(n6173), .C2(n6172), .A(n6171), .B(n6170), .ZN(
        btb_cache_data_in[31]) );
  INV_X1 U4817 ( .A(btb_cache_data_out_rw[30]), .ZN(n6172) );
  INV_X1 U4818 ( .A(n6169), .ZN(n6173) );
  OAI22_X1 U4819 ( .A1(n6445), .A2(n7440), .B1(n4073), .B2(n3942), .ZN(n2642)
         );
  OAI22_X1 U4820 ( .A1(n6464), .A2(n7440), .B1(n4080), .B2(n3942), .ZN(n2650)
         );
  OAI22_X1 U4821 ( .A1(n6451), .A2(n7440), .B1(n4063), .B2(n3942), .ZN(n2645)
         );
  OAI22_X1 U4822 ( .A1(n6436), .A2(n7440), .B1(n4066), .B2(n7439), .ZN(n2639)
         );
  OAI22_X1 U4823 ( .A1(n6454), .A2(n7440), .B1(n6453), .B2(n3938), .ZN(n2646)
         );
  OAI22_X1 U4824 ( .A1(n6460), .A2(n7440), .B1(n6459), .B2(n7439), .ZN(n2648)
         );
  OAI22_X1 U4825 ( .A1(n6449), .A2(n7440), .B1(n4082), .B2(n3938), .ZN(n2644)
         );
  OAI22_X1 U4826 ( .A1(n7106), .A2(n7440), .B1(n4087), .B2(n7439), .ZN(n2651)
         );
  OAI22_X1 U4827 ( .A1(n6434), .A2(n7440), .B1(n4081), .B2(n7439), .ZN(n2638)
         );
  OAI22_X1 U4828 ( .A1(n6428), .A2(n7440), .B1(n4075), .B2(n3938), .ZN(n2634)
         );
  OAI22_X1 U4829 ( .A1(n6430), .A2(n7440), .B1(n4085), .B2(n3942), .ZN(n2635)
         );
  OAI22_X1 U4830 ( .A1(n6439), .A2(n7440), .B1(n4079), .B2(n7439), .ZN(n2640)
         );
  OAI22_X1 U4831 ( .A1(n6457), .A2(n7440), .B1(n6456), .B2(n3942), .ZN(n2647)
         );
  OAI22_X1 U4832 ( .A1(n6469), .A2(n7440), .B1(n4072), .B2(n3938), .ZN(n2652)
         );
  INV_X1 U4833 ( .A(n6470), .ZN(n6469) );
  OAI22_X1 U4834 ( .A1(n6420), .A2(n7440), .B1(n4084), .B2(n7439), .ZN(n2629)
         );
  OAI22_X1 U4835 ( .A1(n6442), .A2(n7440), .B1(n4088), .B2(n7439), .ZN(n2641)
         );
  OAI22_X1 U4836 ( .A1(n6419), .A2(n7440), .B1(n4062), .B2(n7439), .ZN(n2628)
         );
  OAI22_X1 U4837 ( .A1(n6426), .A2(n7440), .B1(n4076), .B2(n3938), .ZN(n2633)
         );
  OAI22_X1 U4838 ( .A1(n6462), .A2(n7440), .B1(n4071), .B2(n7439), .ZN(n2649)
         );
  OAI22_X1 U4839 ( .A1(n6424), .A2(n7440), .B1(n4086), .B2(n3942), .ZN(n2632)
         );
  NAND2_X1 U4840 ( .A1(btb_cache_update_data), .A2(btb_cache_data_out_rw[28]), 
        .ZN(n6131) );
  OAI22_X1 U4841 ( .A1(n6422), .A2(n7440), .B1(n4077), .B2(n3938), .ZN(n2631)
         );
  OAI21_X1 U4842 ( .B1(n5087), .B2(n3870), .A(n6166), .ZN(
        btb_cache_data_in[29]) );
  OAI22_X1 U4843 ( .A1(n6421), .A2(n7440), .B1(n4078), .B2(n3942), .ZN(n2630)
         );
  OAI22_X1 U4844 ( .A1(n7096), .A2(n7095), .B1(n4377), .B2(n7439), .ZN(n2653)
         );
  AOI21_X1 U4845 ( .B1(n7094), .B2(n7093), .A(alu_comp_sel[1]), .ZN(n7095) );
  NAND2_X1 U4846 ( .A1(n7091), .A2(alu_comp_sel[2]), .ZN(n7094) );
  XNOR2_X1 U4847 ( .A(n5051), .B(n4383), .ZN(n7091) );
  OAI211_X1 U4848 ( .C1(n7090), .C2(n7089), .A(n7088), .B(n7087), .ZN(n7096)
         );
  NAND2_X1 U4849 ( .A1(n3920), .A2(n7092), .ZN(n7085) );
  NOR2_X1 U4850 ( .A1(n7092), .A2(alu_comp_sel[2]), .ZN(n7086) );
  NOR2_X1 U4851 ( .A1(n7084), .A2(alu_comp_sel[0]), .ZN(n7090) );
  AOI22_X1 U4852 ( .A1(n5826), .A2(n7107), .B1(btb_cache_update_data), .B2(
        btb_cache_data_out_rw[0]), .ZN(n5827) );
  INV_X1 U4853 ( .A(n6167), .ZN(n5826) );
  OAI22_X1 U4854 ( .A1(n6417), .A2(n7440), .B1(n4064), .B2(n3938), .ZN(n2626)
         );
  INV_X1 U4855 ( .A(btb_cache_data_out_rw[2]), .ZN(n5850) );
  INV_X1 U4856 ( .A(n6431), .ZN(n6430) );
  INV_X1 U4857 ( .A(btb_cache_data_out_rw[16]), .ZN(n5968) );
  INV_X1 U4858 ( .A(n6437), .ZN(n6436) );
  INV_X1 U4859 ( .A(btb_cache_data_out_rw[12]), .ZN(n5941) );
  INV_X1 U4860 ( .A(btb_cache_data_out_rw[7]), .ZN(n5916) );
  INV_X1 U4861 ( .A(n6427), .ZN(n6426) );
  INV_X1 U4862 ( .A(btb_cache_data_out_rw[18]), .ZN(n6002) );
  INV_X1 U4863 ( .A(btb_cache_data_out_rw[21]), .ZN(n6038) );
  INV_X1 U4864 ( .A(btb_cache_data_out_rw[5]), .ZN(n5893) );
  INV_X1 U4865 ( .A(btb_cache_data_out_rw[14]), .ZN(n5953) );
  INV_X1 U4866 ( .A(btb_cache_data_out_rw[27]), .ZN(n6114) );
  INV_X1 U4867 ( .A(btb_cache_data_out_rw[3]), .ZN(n5864) );
  INV_X1 U4868 ( .A(btb_cache_data_out_rw[9]), .ZN(n5924) );
  INV_X1 U4869 ( .A(btb_cache_data_out_rw[13]), .ZN(n5952) );
  INV_X1 U4870 ( .A(btb_cache_data_out_rw[6]), .ZN(n5905) );
  INV_X1 U4871 ( .A(btb_cache_data_out_rw[26]), .ZN(n6112) );
  INV_X1 U4872 ( .A(btb_cache_data_out_rw[1]), .ZN(n5836) );
  INV_X1 U4873 ( .A(n6423), .ZN(n6422) );
  INV_X1 U4874 ( .A(btb_cache_data_out_rw[20]), .ZN(n6028) );
  INV_X1 U4875 ( .A(btb_cache_data_out_rw[24]), .ZN(n6087) );
  INV_X1 U4876 ( .A(btb_cache_data_out_rw[15]), .ZN(n5954) );
  INV_X1 U4877 ( .A(n6443), .ZN(n6442) );
  INV_X1 U4878 ( .A(btb_cache_data_out_rw[10]), .ZN(n5927) );
  INV_X1 U4879 ( .A(btb_cache_data_out_rw[4]), .ZN(n5881) );
  INV_X1 U4880 ( .A(btb_cache_data_out_rw[22]), .ZN(n6054) );
  INV_X1 U4881 ( .A(n6425), .ZN(n6424) );
  INV_X1 U4882 ( .A(btb_cache_data_out_rw[19]), .ZN(n6019) );
  INV_X1 U4883 ( .A(btb_cache_data_out_rw[25]), .ZN(n6097) );
  INV_X1 U4884 ( .A(n6440), .ZN(n6439) );
  INV_X1 U4885 ( .A(btb_cache_data_out_rw[11]), .ZN(n5938) );
  INV_X1 U4886 ( .A(n6429), .ZN(n6428) );
  INV_X1 U4887 ( .A(btb_cache_data_out_rw[17]), .ZN(n5985) );
  INV_X1 U4888 ( .A(btb_cache_data_out_rw[8]), .ZN(n5920) );
  NAND2_X1 U4889 ( .A1(n5044), .A2(btb_cache_update_line), .ZN(n6167) );
  INV_X1 U4890 ( .A(btb_cache_update_line), .ZN(n6171) );
  INV_X1 U4891 ( .A(btb_cache_data_out_rw[23]), .ZN(n6072) );
  OAI22_X1 U4892 ( .A1(n6418), .A2(n7440), .B1(n4065), .B2(n3942), .ZN(n2627)
         );
  OAI22_X1 U4893 ( .A1(n6416), .A2(n7440), .B1(n4067), .B2(n3942), .ZN(n2625)
         );
  OAI22_X1 U4894 ( .A1(n4500), .A2(n7185), .B1(n7184), .B2(n4360), .ZN(n3058)
         );
  OAI22_X1 U4895 ( .A1(n4518), .A2(n7185), .B1(n7184), .B2(n4138), .ZN(n3071)
         );
  OAI22_X1 U4896 ( .A1(n4498), .A2(n7185), .B1(n7184), .B2(n4083), .ZN(n3062)
         );
  OAI22_X1 U4897 ( .A1(n4490), .A2(n7185), .B1(n7184), .B2(n4366), .ZN(n3059)
         );
  OAI22_X1 U4898 ( .A1(n4499), .A2(n7185), .B1(n7184), .B2(n4370), .ZN(n3060)
         );
  OAI22_X1 U4899 ( .A1(n4497), .A2(n7185), .B1(n7184), .B2(n4359), .ZN(n3068)
         );
  OAI22_X1 U4900 ( .A1(n4496), .A2(n7185), .B1(n7184), .B2(n4212), .ZN(n3069)
         );
  OAI22_X1 U4901 ( .A1(n4495), .A2(n7185), .B1(n7184), .B2(n4365), .ZN(n3070)
         );
  OAI22_X1 U4902 ( .A1(n4517), .A2(n7185), .B1(n7184), .B2(n7172), .ZN(n3072)
         );
  OAI22_X1 U4903 ( .A1(n4489), .A2(n7185), .B1(n7184), .B2(n4402), .ZN(n3061)
         );
  NAND2_X1 U4904 ( .A1(n7171), .A2(n4934), .ZN(n7184) );
  NAND2_X1 U4905 ( .A1(n7171), .A2(\ctrl_u/if_stall ), .ZN(n7185) );
  OAI22_X1 U4906 ( .A1(n6476), .A2(n7062), .B1(n4169), .B2(n3942), .ZN(n2818)
         );
  OAI22_X1 U4907 ( .A1(n6409), .A2(n7440), .B1(n4096), .B2(n3942), .ZN(n2622)
         );
  INV_X1 U4908 ( .A(n6410), .ZN(n6409) );
  OAI22_X1 U4909 ( .A1(n6414), .A2(n7440), .B1(n4068), .B2(n3938), .ZN(n2624)
         );
  INV_X1 U4910 ( .A(\dp/pc_plus4_out_if_int[20] ), .ZN(n7129) );
  OAI211_X1 U4911 ( .C1(\intadd_2/SUM[11] ), .C2(n3937), .A(n6377), .B(n6376), 
        .ZN(n2545) );
  AOI22_X1 U4912 ( .A1(n3883), .A2(n6437), .B1(n3928), .B2(
        \dp/pc_plus4_out_if_int[12] ), .ZN(n6376) );
  OAI22_X1 U4913 ( .A1(n3873), .A2(\intadd_2/B[20] ), .B1(\intadd_2/SUM[20] ), 
        .B2(n3879), .ZN(n6400) );
  OAI22_X1 U4914 ( .A1(n5416), .A2(n5393), .B1(\ctrl_u/curr_exe[3] ), .B2(
        n3882), .ZN(\ctrl_u/n458 ) );
  INV_X1 U4915 ( .A(n5392), .ZN(n5393) );
  OAI22_X1 U4916 ( .A1(n5416), .A2(n5391), .B1(\ctrl_u/curr_exe[2] ), .B2(
        n3882), .ZN(\ctrl_u/n459 ) );
  INV_X1 U4917 ( .A(n5390), .ZN(n5391) );
  OAI22_X1 U4918 ( .A1(n5416), .A2(n5406), .B1(cond_sel_exe[1]), .B2(n3882), 
        .ZN(\ctrl_u/n436 ) );
  OAI22_X1 U4919 ( .A1(n5420), .A2(n4126), .B1(n5413), .B2(n4478), .ZN(n5406)
         );
  OAI22_X1 U4920 ( .A1(n5416), .A2(n5398), .B1(\ctrl_u/curr_exe[15] ), .B2(
        n5414), .ZN(\ctrl_u/n446 ) );
  OAI22_X1 U4921 ( .A1(n5420), .A2(n4167), .B1(n5413), .B2(n4454), .ZN(n5398)
         );
  OAI22_X1 U4922 ( .A1(n5416), .A2(n5405), .B1(cond_sel_exe[0]), .B2(n3882), 
        .ZN(\ctrl_u/n437 ) );
  OAI22_X1 U4923 ( .A1(n5420), .A2(n4123), .B1(n5413), .B2(n4491), .ZN(n5405)
         );
  OAI22_X1 U4924 ( .A1(n5416), .A2(n5403), .B1(alu_comp_sel[1]), .B2(n5414), 
        .ZN(\ctrl_u/n439 ) );
  INV_X1 U4925 ( .A(n5402), .ZN(n5403) );
  OAI22_X1 U4926 ( .A1(n5416), .A2(n5395), .B1(\ctrl_u/curr_exe[4] ), .B2(
        n3882), .ZN(\ctrl_u/n457 ) );
  INV_X1 U4927 ( .A(n5394), .ZN(n5395) );
  OAI22_X1 U4928 ( .A1(n5416), .A2(n5397), .B1(\ctrl_u/curr_exe[6] ), .B2(
        n5414), .ZN(\ctrl_u/n455 ) );
  INV_X1 U4929 ( .A(n5396), .ZN(n5397) );
  OAI22_X1 U4930 ( .A1(n5416), .A2(n5415), .B1(shift_type_exe[1]), .B2(n3882), 
        .ZN(\ctrl_u/n426 ) );
  OAI22_X1 U4931 ( .A1(n5420), .A2(n4445), .B1(n5413), .B2(n4522), .ZN(n5415)
         );
  OAI22_X1 U4932 ( .A1(n5416), .A2(n5401), .B1(\ctrl_u/curr_exe[18] ), .B2(
        n5414), .ZN(\ctrl_u/n443 ) );
  INV_X1 U4933 ( .A(n5400), .ZN(n5401) );
  OAI22_X1 U4934 ( .A1(n5416), .A2(n5411), .B1(\ctrl_u/op_type_exe[1] ), .B2(
        n5414), .ZN(\ctrl_u/n432 ) );
  OAI21_X1 U4935 ( .B1(n5420), .B2(op_type_exe[1]), .A(n5410), .ZN(n5411) );
  OAI22_X1 U4936 ( .A1(n5416), .A2(n5399), .B1(\ctrl_u/curr_exe[17] ), .B2(
        n3882), .ZN(\ctrl_u/n444 ) );
  OAI22_X1 U4937 ( .A1(n5420), .A2(n4182), .B1(n5413), .B2(n4484), .ZN(n5399)
         );
  OAI22_X1 U4938 ( .A1(n5416), .A2(n5409), .B1(cond_sel_exe[2]), .B2(n5414), 
        .ZN(\ctrl_u/n435 ) );
  INV_X1 U4939 ( .A(n5408), .ZN(n5409) );
  INV_X1 U4940 ( .A(n5420), .ZN(n5407) );
  OAI22_X1 U4941 ( .A1(n5416), .A2(n5404), .B1(alu_comp_sel[2]), .B2(n3882), 
        .ZN(\ctrl_u/n438 ) );
  OAI22_X1 U4942 ( .A1(n5420), .A2(n4139), .B1(n5413), .B2(n4492), .ZN(n5404)
         );
  OAI22_X1 U4943 ( .A1(n5416), .A2(n5412), .B1(shift_type_exe[0]), .B2(n3882), 
        .ZN(\ctrl_u/n427 ) );
  OAI22_X1 U4944 ( .A1(n5420), .A2(n4378), .B1(n5413), .B2(n4521), .ZN(n5412)
         );
  NOR2_X1 U4945 ( .A1(n5026), .A2(n4867), .ZN(n4922) );
  NAND2_X1 U4946 ( .A1(alu_comp_sel[1]), .A2(alu_comp_sel[2]), .ZN(n7089) );
  AOI22_X1 U4947 ( .A1(n7098), .A2(\dp/a_neg_mult_id_exe_int[18] ), .B1(n7097), 
        .B2(n6431), .ZN(n1458) );
  AOI22_X1 U4948 ( .A1(n7098), .A2(\dp/a_neg_mult_id_exe_int[21] ), .B1(n5194), 
        .B2(n6425), .ZN(n1455) );
  AOI22_X1 U4949 ( .A1(n7098), .A2(\dp/a_neg_mult_id_exe_int[20] ), .B1(n5194), 
        .B2(n6427), .ZN(n1456) );
  AOI22_X1 U4950 ( .A1(n7098), .A2(\dp/a_neg_mult_id_exe_int[16] ), .B1(n7097), 
        .B2(n4891), .ZN(n1460) );
  AOI22_X1 U4951 ( .A1(n7098), .A2(\dp/a_neg_mult_id_exe_int[15] ), .B1(n5194), 
        .B2(n4890), .ZN(n1461) );
  NOR2_X1 U4952 ( .A1(n3937), .A2(\intadd_2/SUM[21] ), .ZN(n5018) );
  XNOR2_X1 U4953 ( .A(n4779), .B(n4778), .ZN(\intadd_2/SUM[21] ) );
  XNOR2_X1 U4954 ( .A(n4356), .B(\dp/imm_id_exe_int[24] ), .ZN(n4778) );
  AOI21_X1 U4955 ( .B1(n4032), .B2(n4824), .A(n4822), .ZN(n4779) );
  NOR2_X1 U4956 ( .A1(n3873), .A2(n4520), .ZN(n5004) );
  NOR2_X1 U4957 ( .A1(\intadd_2/SUM[24] ), .A2(n3879), .ZN(n6401) );
  AOI22_X1 U4958 ( .A1(n5621), .A2(\ctrl_u/next_exe[38] ), .B1(n5622), .B2(
        sub_add_exe), .ZN(\ctrl_u/n423 ) );
  OAI22_X1 U4959 ( .A1(n5132), .A2(n7115), .B1(n366), .B2(n5177), .ZN(n3034)
         );
  INV_X1 U4960 ( .A(\dp/pc_plus4_out_if_int[6] ), .ZN(n7115) );
  OAI22_X1 U4961 ( .A1(n5132), .A2(n7117), .B1(n368), .B2(n5177), .ZN(n3032)
         );
  INV_X1 U4962 ( .A(\dp/pc_plus4_out_if_int[8] ), .ZN(n7117) );
  OAI22_X1 U4963 ( .A1(n5131), .A2(n7110), .B1(n361), .B2(n5177), .ZN(n3039)
         );
  INV_X1 U4964 ( .A(\dp/pc_plus4_out_if_int[1] ), .ZN(n7110) );
  OAI22_X1 U4965 ( .A1(n5132), .A2(btb_cache_read_address[0]), .B1(n360), .B2(
        n5177), .ZN(n3040) );
  OAI22_X1 U4966 ( .A1(n5131), .A2(n7112), .B1(n363), .B2(n5177), .ZN(n3037)
         );
  INV_X1 U4967 ( .A(\dp/pc_plus4_out_if_int[3] ), .ZN(n7112) );
  OAI22_X1 U4968 ( .A1(n5131), .A2(n7116), .B1(n367), .B2(n5177), .ZN(n3033)
         );
  INV_X1 U4969 ( .A(\dp/pc_plus4_out_if_int[7] ), .ZN(n7116) );
  OAI22_X1 U4970 ( .A1(n5132), .A2(n7113), .B1(n364), .B2(n5177), .ZN(n3036)
         );
  INV_X1 U4971 ( .A(\dp/pc_plus4_out_if_int[4] ), .ZN(n7113) );
  OAI22_X1 U4972 ( .A1(n5130), .A2(n7111), .B1(n362), .B2(n5177), .ZN(n3038)
         );
  INV_X1 U4973 ( .A(\dp/pc_plus4_out_if_int[2] ), .ZN(n7111) );
  OAI22_X1 U4974 ( .A1(n5131), .A2(n7114), .B1(n365), .B2(n5177), .ZN(n3035)
         );
  INV_X1 U4975 ( .A(\dp/pc_plus4_out_if_int[5] ), .ZN(n7114) );
  INV_X1 U4976 ( .A(n7182), .ZN(n281) );
  AOI22_X1 U4977 ( .A1(n5133), .A2(rs_id[2]), .B1(n5180), .B2(instr_if[23]), 
        .ZN(n7182) );
  AOI22_X1 U4978 ( .A1(n5621), .A2(\ctrl_u/next_exe[5] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[5] ), .ZN(\ctrl_u/n456 ) );
  AOI22_X1 U4979 ( .A1(n5621), .A2(\ctrl_u/next_exe[1] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[1] ), .ZN(\ctrl_u/n460 ) );
  AOI22_X1 U4980 ( .A1(n5621), .A2(\ctrl_u/next_exe[0] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[0] ), .ZN(\ctrl_u/n461 ) );
  AOI22_X1 U4981 ( .A1(n5621), .A2(\ctrl_u/next_exe[36] ), .B1(n5622), .B2(
        shift_type_exe[2]), .ZN(\ctrl_u/n425 ) );
  OAI211_X1 U4982 ( .C1(\intadd_2/SUM[9] ), .C2(n3937), .A(n6373), .B(n6372), 
        .ZN(n2547) );
  AOI22_X1 U4983 ( .A1(n3883), .A2(n6443), .B1(n3936), .B2(
        \dp/pc_plus4_out_if_int[10] ), .ZN(n6372) );
  OAI211_X1 U4984 ( .C1(\intadd_2/SUM[10] ), .C2(n3937), .A(n6375), .B(n6374), 
        .ZN(n2546) );
  AOI22_X1 U4985 ( .A1(n3883), .A2(n6440), .B1(n3936), .B2(
        \dp/pc_plus4_out_if_int[11] ), .ZN(n6374) );
  OAI211_X1 U4986 ( .C1(\intadd_2/SUM[16] ), .C2(n3937), .A(n6392), .B(n6391), 
        .ZN(n2540) );
  AOI22_X1 U4987 ( .A1(n3883), .A2(n6429), .B1(n3928), .B2(
        \dp/pc_plus4_out_if_int[17] ), .ZN(n6391) );
  OAI21_X1 U4988 ( .B1(n5984), .B2(n6027), .A(n5983), .ZN(n6429) );
  AOI21_X1 U4989 ( .B1(n3954), .B2(\dp/exs/alu_unit/shifter_out[19] ), .A(
        n5982), .ZN(n5983) );
  OAI21_X1 U4990 ( .B1(\intadd_1/SUM[18] ), .B2(n7066), .A(n5981), .ZN(n5982)
         );
  NAND2_X1 U4991 ( .A1(n5978), .A2(n3952), .ZN(n5979) );
  AOI211_X1 U4992 ( .C1(\dp/exs/alu_unit/shifter_out[0] ), .C2(n3954), .A(
        n7082), .B(n7081), .ZN(n7084) );
  OAI211_X1 U4993 ( .C1(n7080), .C2(n7079), .A(n7078), .B(n7077), .ZN(n7081)
         );
  NAND2_X1 U4994 ( .A1(n7076), .A2(n7075), .ZN(n7077) );
  OAI21_X1 U4995 ( .B1(n4369), .B2(n5169), .A(n7074), .ZN(n7075) );
  OAI21_X1 U4996 ( .B1(\dp/b10_1_mult_id_exe_int[1] ), .B2(n5150), .A(n7073), 
        .ZN(n7074) );
  NAND2_X1 U4997 ( .A1(n7070), .A2(n3953), .ZN(n7078) );
  OAI22_X1 U4998 ( .A1(n7070), .A2(n7068), .B1(n7067), .B2(n7066), .ZN(n7082)
         );
  NAND2_X1 U4999 ( .A1(n7071), .A2(n3952), .ZN(n7068) );
  INV_X1 U5000 ( .A(n7079), .ZN(n7065) );
  AOI21_X1 U5001 ( .B1(n5621), .B2(n6327), .A(n5344), .ZN(n5345) );
  OAI22_X1 U5002 ( .A1(n5130), .A2(n3854), .B1(n389), .B2(n5177), .ZN(n3011)
         );
  OAI22_X1 U5003 ( .A1(n5132), .A2(n7173), .B1(n5177), .B2(n7172), .ZN(n274)
         );
  INV_X1 U5004 ( .A(instr_if[16]), .ZN(n7173) );
  OAI22_X1 U5005 ( .A1(n5131), .A2(n7175), .B1(n5177), .B2(n4365), .ZN(n276)
         );
  INV_X1 U5006 ( .A(instr_if[18]), .ZN(n7175) );
  OAI22_X1 U5007 ( .A1(n5131), .A2(n7174), .B1(n5177), .B2(n4138), .ZN(n275)
         );
  INV_X1 U5008 ( .A(instr_if[17]), .ZN(n7174) );
  NAND2_X1 U5009 ( .A1(n4057), .A2(n6754), .ZN(n2884) );
  NAND2_X1 U5010 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[62] ), .ZN(n6754) );
  NAND2_X1 U5011 ( .A1(n4057), .A2(n6724), .ZN(n2914) );
  NAND2_X1 U5012 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[32] ), .ZN(n6724) );
  OAI22_X1 U5013 ( .A1(n5131), .A2(n7133), .B1(n384), .B2(n5177), .ZN(n3016)
         );
  INV_X1 U5014 ( .A(\dp/pc_plus4_out_if_int[24] ), .ZN(n7133) );
  OAI22_X1 U5015 ( .A1(n5131), .A2(n7134), .B1(n385), .B2(n5178), .ZN(n3015)
         );
  INV_X1 U5016 ( .A(\dp/pc_plus4_out_if_int[25] ), .ZN(n7134) );
  OAI22_X1 U5017 ( .A1(n5132), .A2(n7136), .B1(n387), .B2(n5177), .ZN(n3013)
         );
  INV_X1 U5018 ( .A(\dp/pc_plus4_out_if_int[27] ), .ZN(n7136) );
  OAI22_X1 U5019 ( .A1(n5132), .A2(n7135), .B1(n386), .B2(n5177), .ZN(n3014)
         );
  INV_X1 U5020 ( .A(\dp/pc_plus4_out_if_int[26] ), .ZN(n7135) );
  OAI22_X1 U5021 ( .A1(n5131), .A2(n7132), .B1(n383), .B2(n4850), .ZN(n3017)
         );
  INV_X1 U5022 ( .A(\dp/pc_plus4_out_if_int[23] ), .ZN(n7132) );
  OAI22_X1 U5023 ( .A1(n5132), .A2(n7131), .B1(n382), .B2(n4850), .ZN(n3018)
         );
  INV_X1 U5024 ( .A(\dp/pc_plus4_out_if_int[22] ), .ZN(n7131) );
  OAI22_X1 U5025 ( .A1(n5130), .A2(n7137), .B1(n388), .B2(n5177), .ZN(n3012)
         );
  INV_X1 U5026 ( .A(\dp/pc_plus4_out_if_int[28] ), .ZN(n7137) );
  OAI21_X1 U5027 ( .B1(n3934), .B2(n4502), .A(n5539), .ZN(\ctrl_u/n508 ) );
  OAI22_X1 U5028 ( .A1(n5132), .A2(n7176), .B1(n4212), .B2(n5177), .ZN(n277)
         );
  INV_X1 U5029 ( .A(instr_if[19]), .ZN(n7176) );
  OAI22_X1 U5030 ( .A1(n5131), .A2(n7178), .B1(n4651), .B2(n4359), .ZN(n278)
         );
  INV_X1 U5031 ( .A(instr_if[20]), .ZN(n7178) );
  OAI22_X1 U5032 ( .A1(n5132), .A2(n7125), .B1(n376), .B2(n5177), .ZN(n3024)
         );
  INV_X1 U5033 ( .A(\dp/pc_plus4_out_if_int[16] ), .ZN(n7125) );
  OAI22_X1 U5034 ( .A1(n5132), .A2(n7119), .B1(n370), .B2(n4850), .ZN(n3030)
         );
  INV_X1 U5035 ( .A(\dp/pc_plus4_out_if_int[10] ), .ZN(n7119) );
  OAI22_X1 U5036 ( .A1(n5131), .A2(n7118), .B1(n369), .B2(n5177), .ZN(n3031)
         );
  INV_X1 U5037 ( .A(\dp/pc_plus4_out_if_int[9] ), .ZN(n7118) );
  OAI22_X1 U5038 ( .A1(n5132), .A2(n7120), .B1(n371), .B2(n4850), .ZN(n3029)
         );
  INV_X1 U5039 ( .A(\dp/pc_plus4_out_if_int[11] ), .ZN(n7120) );
  OAI22_X1 U5040 ( .A1(n5131), .A2(n7121), .B1(n372), .B2(n4850), .ZN(n3028)
         );
  INV_X1 U5041 ( .A(\dp/pc_plus4_out_if_int[12] ), .ZN(n7121) );
  OAI22_X1 U5042 ( .A1(n5131), .A2(n7130), .B1(n381), .B2(n4850), .ZN(n3019)
         );
  INV_X1 U5043 ( .A(\dp/pc_plus4_out_if_int[21] ), .ZN(n7130) );
  OAI22_X1 U5044 ( .A1(n5132), .A2(n7127), .B1(n378), .B2(n5177), .ZN(n3022)
         );
  INV_X1 U5045 ( .A(\dp/pc_plus4_out_if_int[18] ), .ZN(n7127) );
  OAI22_X1 U5046 ( .A1(n5131), .A2(n7122), .B1(n373), .B2(n5177), .ZN(n3027)
         );
  INV_X1 U5047 ( .A(\dp/pc_plus4_out_if_int[13] ), .ZN(n7122) );
  OAI22_X1 U5048 ( .A1(n5131), .A2(n7128), .B1(n379), .B2(n5177), .ZN(n3021)
         );
  INV_X1 U5049 ( .A(\dp/pc_plus4_out_if_int[19] ), .ZN(n7128) );
  OAI22_X1 U5050 ( .A1(n5131), .A2(n7124), .B1(n375), .B2(n5177), .ZN(n3025)
         );
  INV_X1 U5051 ( .A(\dp/pc_plus4_out_if_int[15] ), .ZN(n7124) );
  OAI22_X1 U5052 ( .A1(n5132), .A2(n7123), .B1(n374), .B2(n4651), .ZN(n3026)
         );
  INV_X1 U5053 ( .A(\dp/pc_plus4_out_if_int[14] ), .ZN(n7123) );
  OAI22_X1 U5054 ( .A1(n5132), .A2(n7126), .B1(n377), .B2(n5177), .ZN(n3023)
         );
  INV_X1 U5055 ( .A(\dp/pc_plus4_out_if_int[17] ), .ZN(n7126) );
  NAND2_X1 U5056 ( .A1(n6786), .A2(n6785), .ZN(n2920) );
  NAND2_X1 U5057 ( .A1(n5202), .A2(n6784), .ZN(n6785) );
  INV_X1 U5058 ( .A(n6788), .ZN(n6784) );
  NAND2_X1 U5059 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[26] ), .ZN(n6786) );
  NAND2_X1 U5060 ( .A1(n6819), .A2(n6818), .ZN(n2926) );
  NAND2_X1 U5061 ( .A1(n5202), .A2(n6817), .ZN(n6818) );
  INV_X1 U5062 ( .A(n6821), .ZN(n6817) );
  NAND2_X1 U5063 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[20] ), .ZN(n6819) );
  AOI22_X1 U5064 ( .A1(n5126), .A2(\dp/a_neg_mult_id_exe_int[22] ), .B1(n5194), 
        .B2(n6423), .ZN(n1454) );
  AOI22_X1 U5065 ( .A1(n5126), .A2(\dp/a_neg_mult_id_exe_int[1] ), .B1(n5194), 
        .B2(n6470), .ZN(n1475) );
  NAND2_X1 U5066 ( .A1(n5473), .A2(n4815), .ZN(\ctrl_u/n533 ) );
  NOR3_X1 U5067 ( .A1(n5637), .A2(n5471), .A3(n5470), .ZN(n5472) );
  OAI21_X1 U5068 ( .B1(n5504), .B2(n7275), .A(n5469), .ZN(n5470) );
  AOI211_X1 U5069 ( .C1(n5504), .C2(n5590), .A(n5553), .B(n5647), .ZN(n5469)
         );
  AOI21_X1 U5070 ( .B1(n5498), .B2(n5468), .A(n5594), .ZN(n5471) );
  INV_X1 U5071 ( .A(n5467), .ZN(n5468) );
  NAND2_X1 U5072 ( .A1(n5479), .A2(n4815), .ZN(\ctrl_u/n530 ) );
  NOR3_X1 U5073 ( .A1(n5637), .A2(n5477), .A3(n5476), .ZN(n5478) );
  NOR2_X1 U5074 ( .A1(n7289), .A2(n5594), .ZN(n5477) );
  NAND2_X1 U5075 ( .A1(n5454), .A2(n4815), .ZN(\ctrl_u/n534 ) );
  AOI211_X1 U5076 ( .C1(n5499), .C2(n5452), .A(n5637), .B(n5451), .ZN(n5453)
         );
  OAI211_X1 U5077 ( .C1(instr_if[16]), .C2(n5450), .A(n5635), .B(n5449), .ZN(
        n5451) );
  AOI211_X1 U5078 ( .C1(n5649), .C2(instr_if[28]), .A(n5448), .B(n5447), .ZN(
        n5449) );
  NOR2_X1 U5079 ( .A1(instr_if[28]), .A2(n5644), .ZN(n5447) );
  AOI21_X1 U5080 ( .B1(n5627), .B2(n5446), .A(n5590), .ZN(n5448) );
  INV_X1 U5081 ( .A(n5588), .ZN(n5446) );
  OR4_X1 U5082 ( .A1(instr_if[1]), .A2(n7295), .A3(n5455), .A4(n5444), .ZN(
        n5452) );
  INV_X1 U5083 ( .A(n5585), .ZN(n5444) );
  NAND2_X1 U5084 ( .A1(n5426), .A2(n5425), .ZN(\ctrl_u/n510 ) );
  INV_X1 U5085 ( .A(n5525), .ZN(n5424) );
  OAI21_X1 U5086 ( .B1(n5599), .B2(n4448), .A(n5425), .ZN(\ctrl_u/n509 ) );
  NOR2_X1 U5087 ( .A1(n5619), .A2(n5423), .ZN(n5425) );
  NOR3_X1 U5088 ( .A1(n5422), .A2(n5481), .A3(\ctrl_u/if_stall ), .ZN(n5423)
         );
  OAI211_X1 U5089 ( .C1(\intadd_2/SUM[17] ), .C2(n3937), .A(n6394), .B(n6393), 
        .ZN(n2539) );
  AOI22_X1 U5090 ( .A1(n3884), .A2(n6427), .B1(n3928), .B2(
        \dp/pc_plus4_out_if_int[18] ), .ZN(n6393) );
  OAI21_X1 U5091 ( .B1(n6001), .B2(n6027), .A(n6000), .ZN(n6427) );
  AOI21_X1 U5092 ( .B1(n3954), .B2(\dp/exs/alu_unit/shifter_out[20] ), .A(
        n5999), .ZN(n6000) );
  OAI21_X1 U5093 ( .B1(\intadd_1/SUM[19] ), .B2(n7066), .A(n5998), .ZN(n5999)
         );
  NAND2_X1 U5094 ( .A1(n5995), .A2(n3952), .ZN(n5996) );
  NAND2_X1 U5095 ( .A1(n4903), .A2(n5006), .ZN(n6003) );
  NAND2_X1 U5096 ( .A1(n5988), .A2(n5007), .ZN(n4903) );
  OAI211_X1 U5097 ( .C1(\intadd_2/SUM[15] ), .C2(n3937), .A(n6390), .B(n6389), 
        .ZN(n2541) );
  AOI22_X1 U5098 ( .A1(n3883), .A2(n6431), .B1(n3936), .B2(
        \dp/pc_plus4_out_if_int[16] ), .ZN(n6389) );
  OAI21_X1 U5099 ( .B1(n5967), .B2(n6027), .A(n5966), .ZN(n6431) );
  AOI21_X1 U5100 ( .B1(\dp/exs/alu_unit/shifter_out[18] ), .B2(n7083), .A(
        n5965), .ZN(n5966) );
  OAI21_X1 U5101 ( .B1(n3862), .B2(n7066), .A(n5964), .ZN(n5965) );
  NAND2_X1 U5102 ( .A1(n5961), .A2(n3952), .ZN(n5962) );
  AOI22_X1 U5103 ( .A1(n5647), .A2(n5516), .B1(n5534), .B2(n5515), .ZN(n5517)
         );
  NOR2_X1 U5104 ( .A1(instr_if[3]), .A2(n7281), .ZN(n5515) );
  NOR2_X1 U5105 ( .A1(n5514), .A2(n5543), .ZN(n5516) );
  AOI22_X1 U5106 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[5] ), .B1(n5194), 
        .B2(n4883), .ZN(n1471) );
  AOI22_X1 U5107 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[14] ), .B1(n7097), 
        .B2(n6437), .ZN(n1462) );
  AOI22_X1 U5108 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[13] ), .B1(n5194), 
        .B2(n6440), .ZN(n1463) );
  OAI21_X1 U5109 ( .B1(n5937), .B2(n6027), .A(n5936), .ZN(n6440) );
  AOI21_X1 U5110 ( .B1(\dp/exs/alu_unit/shifter_out[13] ), .B2(n3954), .A(
        n5935), .ZN(n5936) );
  OAI21_X1 U5111 ( .B1(\intadd_1/SUM[12] ), .B2(n7066), .A(n5934), .ZN(n5935)
         );
  NAND2_X1 U5112 ( .A1(n4936), .A2(n3952), .ZN(n5932) );
  INV_X1 U5113 ( .A(n4935), .ZN(n4936) );
  OAI21_X1 U5114 ( .B1(n4935), .B2(n3953), .A(n4937), .ZN(n5933) );
  NAND2_X1 U5115 ( .A1(n4935), .A2(n7080), .ZN(n4937) );
  BUF_X1 U5116 ( .A(n4938), .Z(n4935) );
  AOI22_X1 U5117 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[12] ), .B1(n5194), 
        .B2(n6443), .ZN(n1464) );
  AOI22_X1 U5118 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[2] ), .B1(n7097), 
        .B2(n4892), .ZN(n1474) );
  AOI22_X1 U5119 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[3] ), .B1(n5194), 
        .B2(n4881), .ZN(n1473) );
  AOI22_X1 U5120 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[4] ), .B1(n5194), 
        .B2(n4882), .ZN(n1472) );
  AOI22_X1 U5121 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[11] ), .B1(n5194), 
        .B2(n4889), .ZN(n1465) );
  AOI22_X1 U5122 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[8] ), .B1(n5194), 
        .B2(n4886), .ZN(n1468) );
  AOI22_X1 U5123 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[9] ), .B1(n5194), 
        .B2(n4887), .ZN(n1467) );
  AOI22_X1 U5124 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[6] ), .B1(n5194), 
        .B2(n4884), .ZN(n1470) );
  AOI22_X1 U5125 ( .A1(n5127), .A2(\dp/a_neg_mult_id_exe_int[7] ), .B1(n5194), 
        .B2(n4885), .ZN(n1469) );
  AOI22_X1 U5126 ( .A1(\dp/a_neg_mult_id_exe_int[23] ), .A2(n5126), .B1(n4900), 
        .B2(n5194), .ZN(n1453) );
  OAI21_X1 U5127 ( .B1(n6979), .B2(n5204), .A(n6978), .ZN(n2660) );
  NAND2_X1 U5128 ( .A1(n5209), .A2(\dp/b_adder_id_exe_int[25] ), .ZN(n6978) );
  OAI21_X1 U5129 ( .B1(n7042), .B2(n5203), .A(n7041), .ZN(n2681) );
  NAND2_X1 U5130 ( .A1(n5210), .A2(\dp/b_adder_id_exe_int[4] ), .ZN(n7041) );
  OAI21_X1 U5131 ( .B1(n6844), .B2(n5204), .A(n6843), .ZN(n2868) );
  NAND2_X1 U5132 ( .A1(n5210), .A2(n4250), .ZN(n6843) );
  OAI21_X1 U5133 ( .B1(n6841), .B2(n5205), .A(n6840), .ZN(n2867) );
  NAND2_X1 U5134 ( .A1(n5209), .A2(n4462), .ZN(n6840) );
  AND2_X1 U5135 ( .A1(n5568), .A2(n5567), .ZN(n5569) );
  OAI21_X1 U5136 ( .B1(n6868), .B2(n3875), .A(n6867), .ZN(n2876) );
  NAND2_X1 U5137 ( .A1(n5210), .A2(n4254), .ZN(n6867) );
  OAI21_X1 U5138 ( .B1(n6873), .B2(n3874), .A(n6872), .ZN(n2877) );
  NAND2_X1 U5139 ( .A1(n5209), .A2(n4285), .ZN(n6872) );
  OAI21_X1 U5140 ( .B1(n6847), .B2(n3875), .A(n6846), .ZN(n2869) );
  NAND2_X1 U5141 ( .A1(n5209), .A2(n4251), .ZN(n6846) );
  OAI21_X1 U5142 ( .B1(n6806), .B2(n5203), .A(n6805), .ZN(n2859) );
  NAND2_X1 U5143 ( .A1(n5210), .A2(n4244), .ZN(n6805) );
  OAI21_X1 U5144 ( .B1(n6862), .B2(n5204), .A(n6861), .ZN(n2875) );
  NAND2_X1 U5145 ( .A1(n5209), .A2(n4253), .ZN(n6861) );
  OAI21_X1 U5146 ( .B1(n6782), .B2(n3874), .A(n6781), .ZN(n2855) );
  NAND2_X1 U5147 ( .A1(n5210), .A2(n4459), .ZN(n6781) );
  OAI21_X1 U5148 ( .B1(n6838), .B2(n3875), .A(n6837), .ZN(n2866) );
  NAND2_X1 U5149 ( .A1(n5210), .A2(n4461), .ZN(n6837) );
  OAI21_X1 U5150 ( .B1(n6835), .B2(n5203), .A(n6834), .ZN(n2865) );
  NAND2_X1 U5151 ( .A1(n5209), .A2(n4460), .ZN(n6834) );
  OAI21_X1 U5152 ( .B1(n6800), .B2(n5204), .A(n6799), .ZN(n2858) );
  NAND2_X1 U5153 ( .A1(n5210), .A2(n4243), .ZN(n6799) );
  OAI21_X1 U5154 ( .B1(n6794), .B2(n5205), .A(n6793), .ZN(n2857) );
  NAND2_X1 U5155 ( .A1(n5209), .A2(n4242), .ZN(n6793) );
  AOI22_X1 U5156 ( .A1(\ctrl_u/curr_exe_41 ), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/next_exe[41] ), .ZN(\ctrl_u/n420 ) );
  AOI22_X1 U5157 ( .A1(log_type_exe[3]), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/next_exe[33] ), .ZN(\ctrl_u/n428 ) );
  AOI22_X1 U5158 ( .A1(\ctrl_u/curr_exe_39 ), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/next_exe[39] ), .ZN(\ctrl_u/n422 ) );
  AOI22_X1 U5159 ( .A1(\ctrl_u/curr_ak_exe ), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/curr_ak_id ), .ZN(\ctrl_u/n169 ) );
  AOI22_X1 U5160 ( .A1(log_type_exe[1]), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/next_exe[31] ), .ZN(\ctrl_u/n430 ) );
  AOI22_X1 U5161 ( .A1(\ctrl_u/curr_pt_exe ), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/curr_pt_id ), .ZN(\ctrl_u/n166 ) );
  AOI22_X1 U5162 ( .A1(\ctrl_u/curr_exe_40 ), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/next_exe[40] ), .ZN(\ctrl_u/n421 ) );
  AOI22_X1 U5163 ( .A1(log_type_exe[2]), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/next_exe[32] ), .ZN(\ctrl_u/n429 ) );
  AOI22_X1 U5164 ( .A1(\ctrl_u/curr_exe[19] ), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/next_exe[19] ), .ZN(\ctrl_u/n442 ) );
  AOI22_X1 U5165 ( .A1(op_type_exe[0]), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/next_exe[28] ), .ZN(\ctrl_u/n433 ) );
  AOI21_X1 U5166 ( .B1(\ctrl_u/curr_id[13] ), .B2(n3941), .A(n5551), .ZN(
        \ctrl_u/n386 ) );
  INV_X1 U5167 ( .A(n5557), .ZN(n5551) );
  OAI22_X1 U5168 ( .A1(n5547), .A2(n7281), .B1(n5182), .B2(n4584), .ZN(
        \ctrl_u/n511 ) );
  OAI21_X1 U5169 ( .B1(n7163), .B2(n4398), .A(n7149), .ZN(n3046) );
  OAI22_X1 U5170 ( .A1(n6500), .A2(n7062), .B1(n4171), .B2(n3938), .ZN(n2814)
         );
  OAI22_X1 U5171 ( .A1(n6495), .A2(n7062), .B1(n4170), .B2(n3942), .ZN(n2815)
         );
  NAND2_X1 U5172 ( .A1(n5213), .A2(\dp/ids/rp2[19] ), .ZN(n6915) );
  AOI22_X1 U5173 ( .A1(n3898), .A2(\dp/id_exe_regs/b_mult_reg/q[18] ), .B1(
        n3956), .B2(\dp/id_exe_regs/b_mult_reg/q[20] ), .ZN(n6914) );
  AOI21_X1 U5174 ( .B1(\ctrl_u/curr_id[31] ), .B2(n3941), .A(n5527), .ZN(
        \ctrl_u/n305 ) );
  AOI21_X1 U5175 ( .B1(\ctrl_u/curr_id[32] ), .B2(n3941), .A(n5527), .ZN(
        \ctrl_u/n303 ) );
  AOI222_X1 U5176 ( .A1(n5525), .A2(n5529), .B1(instr_if[0]), .B2(n5524), .C1(
        n5596), .C2(n5523), .ZN(n5526) );
  INV_X1 U5177 ( .A(n5531), .ZN(n5523) );
  NAND2_X1 U5178 ( .A1(n5562), .A2(n5589), .ZN(n5525) );
  OAI22_X1 U5179 ( .A1(n5196), .A2(n6500), .B1(n4472), .B2(n4808), .ZN(n2846)
         );
  XNOR2_X1 U5180 ( .A(n6499), .B(n6498), .ZN(n6500) );
  NAND2_X1 U5181 ( .A1(n6504), .A2(n6497), .ZN(n6498) );
  INV_X1 U5182 ( .A(n6514), .ZN(n6496) );
  AOI21_X1 U5183 ( .B1(\ctrl_u/curr_id[33] ), .B2(n3941), .A(n5528), .ZN(
        \ctrl_u/n301 ) );
  OAI211_X1 U5184 ( .C1(n3935), .C2(n4581), .A(n5539), .B(n5538), .ZN(
        \ctrl_u/n532 ) );
  OR2_X1 U5185 ( .A1(n3927), .A2(n4605), .ZN(n5538) );
  OAI22_X1 U5186 ( .A1(instr_if[2]), .A2(instr_if[0]), .B1(n5596), .B2(n7279), 
        .ZN(n5537) );
  OAI211_X1 U5187 ( .C1(n5649), .C2(n5511), .A(n5651), .B(n5512), .ZN(n5492)
         );
  OAI211_X1 U5188 ( .C1(n5491), .C2(n5506), .A(n5505), .B(n5567), .ZN(n5493)
         );
  AOI22_X1 U5189 ( .A1(n3955), .A2(\dp/ids/rp2[0] ), .B1(n7100), .B2(
        \dp/op_b_id_ex_int[0] ), .ZN(n1144) );
  AOI22_X1 U5190 ( .A1(n3955), .A2(\dp/ids/rp2[1] ), .B1(n7100), .B2(
        \dp/op_b_id_ex_int[1] ), .ZN(n1143) );
  OAI22_X1 U5191 ( .A1(n5563), .A2(n5562), .B1(n5182), .B2(n4543), .ZN(
        \ctrl_u/n548 ) );
  INV_X1 U5192 ( .A(n6590), .ZN(n6592) );
  OAI21_X1 U5193 ( .B1(n6758), .B2(n3874), .A(n6757), .ZN(n2851) );
  NAND2_X1 U5194 ( .A1(n5207), .A2(n4455), .ZN(n6757) );
  AOI22_X1 U5195 ( .A1(n6415), .A2(n5194), .B1(\dp/a_neg_mult_id_exe_int[29] ), 
        .B2(n5126), .ZN(n1447) );
  INV_X1 U5196 ( .A(n6414), .ZN(n6415) );
  AOI22_X1 U5197 ( .A1(n4899), .A2(n5194), .B1(\dp/a_neg_mult_id_exe_int[28] ), 
        .B2(n5126), .ZN(n1448) );
  AOI22_X1 U5198 ( .A1(n4901), .A2(n5194), .B1(\dp/a_neg_mult_id_exe_int[27] ), 
        .B2(n5126), .ZN(n1449) );
  AOI22_X1 U5199 ( .A1(n4893), .A2(n7097), .B1(\dp/a_neg_mult_id_exe_int[24] ), 
        .B2(n5126), .ZN(n1452) );
  OAI211_X1 U5200 ( .C1(\intadd_1/SUM[23] ), .C2(n7066), .A(n6051), .B(n6050), 
        .ZN(n6052) );
  NAND2_X1 U5201 ( .A1(n6047), .A2(n3952), .ZN(n6048) );
  NAND2_X1 U5202 ( .A1(\dp/exs/alu_unit/shifter_out[24] ), .A2(n3954), .ZN(
        n6051) );
  XNOR2_X1 U5203 ( .A(n6056), .B(n6057), .ZN(n6046) );
  AOI22_X1 U5204 ( .A1(n4897), .A2(n5194), .B1(\dp/a_neg_mult_id_exe_int[26] ), 
        .B2(n5126), .ZN(n1450) );
  OAI21_X1 U5205 ( .B1(n5224), .B2(n4399), .A(n7149), .ZN(n3045) );
  OAI21_X1 U5206 ( .B1(n5224), .B2(n4367), .A(n7149), .ZN(n3043) );
  OAI21_X1 U5207 ( .B1(n5225), .B2(n4397), .A(n7149), .ZN(n3047) );
  OAI21_X1 U5208 ( .B1(n5225), .B2(n4503), .A(n7149), .ZN(n3042) );
  OAI21_X1 U5209 ( .B1(n5225), .B2(n4400), .A(n7149), .ZN(n3044) );
  INV_X1 U5210 ( .A(n7147), .ZN(n7148) );
  OAI21_X1 U5211 ( .B1(n6996), .B2(n5205), .A(n6995), .ZN(n2668) );
  NAND2_X1 U5212 ( .A1(n5207), .A2(\dp/b_adder_id_exe_int[17] ), .ZN(n6995) );
  OAI21_X1 U5213 ( .B1(n7001), .B2(n3875), .A(n7000), .ZN(n2669) );
  NAND2_X1 U5214 ( .A1(n5206), .A2(\dp/b_adder_id_exe_int[16] ), .ZN(n7000) );
  OAI22_X1 U5215 ( .A1(n6689), .A2(n7062), .B1(n4178), .B2(n3942), .ZN(n2792)
         );
  OAI22_X1 U5216 ( .A1(n7163), .A2(\intadd_2/A[4] ), .B1(n4375), .B2(n4865), 
        .ZN(n257) );
  OAI22_X1 U5217 ( .A1(n7163), .A2(n4099), .B1(n4376), .B2(n4865), .ZN(n256)
         );
  OAI22_X1 U5218 ( .A1(n7163), .A2(n4070), .B1(n4368), .B2(n4865), .ZN(n265)
         );
  OAI22_X1 U5219 ( .A1(n7163), .A2(\intadd_2/A[6] ), .B1(n4373), .B2(n4865), 
        .ZN(n259) );
  OAI21_X1 U5220 ( .B1(n6770), .B2(n5205), .A(n6769), .ZN(n2853) );
  NAND2_X1 U5221 ( .A1(n5207), .A2(n4457), .ZN(n6769) );
  OAI21_X1 U5222 ( .B1(n6764), .B2(n5203), .A(n6763), .ZN(n2852) );
  NAND2_X1 U5223 ( .A1(n5206), .A2(n4456), .ZN(n6763) );
  OAI21_X1 U5224 ( .B1(n6816), .B2(n3874), .A(n6815), .ZN(n2861) );
  NAND2_X1 U5225 ( .A1(n5207), .A2(n4246), .ZN(n6815) );
  OAI21_X1 U5226 ( .B1(n6811), .B2(n5204), .A(n6810), .ZN(n2860) );
  NAND2_X1 U5227 ( .A1(n5206), .A2(n4245), .ZN(n6810) );
  OAI21_X1 U5228 ( .B1(n6776), .B2(n5205), .A(n6775), .ZN(n2854) );
  NAND2_X1 U5229 ( .A1(n5208), .A2(n4458), .ZN(n6775) );
  OAI21_X1 U5230 ( .B1(n6879), .B2(n3874), .A(n6878), .ZN(n2878) );
  NAND2_X1 U5231 ( .A1(n5206), .A2(n4467), .ZN(n6878) );
  OAI21_X1 U5232 ( .B1(n6821), .B2(n3875), .A(n6820), .ZN(n2862) );
  NAND2_X1 U5233 ( .A1(n5208), .A2(n4247), .ZN(n6820) );
  OAI21_X1 U5234 ( .B1(n6849), .B2(n5203), .A(n6848), .ZN(n2870) );
  NAND2_X1 U5235 ( .A1(n5206), .A2(n4252), .ZN(n6848) );
  OAI21_X1 U5236 ( .B1(n6826), .B2(n3874), .A(n6825), .ZN(n2863) );
  NAND2_X1 U5237 ( .A1(n5207), .A2(n4248), .ZN(n6825) );
  OAI21_X1 U5238 ( .B1(n6884), .B2(n3875), .A(n6883), .ZN(n2880) );
  NAND2_X1 U5239 ( .A1(n5208), .A2(n4469), .ZN(n6883) );
  OAI21_X1 U5240 ( .B1(n6882), .B2(n5203), .A(n6881), .ZN(n2879) );
  NAND2_X1 U5241 ( .A1(n5207), .A2(n4468), .ZN(n6881) );
  OAI21_X1 U5242 ( .B1(n7054), .B2(n5204), .A(n7053), .ZN(n2684) );
  NAND2_X1 U5243 ( .A1(n5207), .A2(\dp/b_adder_id_exe_int[1] ), .ZN(n7053) );
  OAI21_X1 U5244 ( .B1(n6855), .B2(n5205), .A(n6854), .ZN(n2873) );
  NAND2_X1 U5245 ( .A1(n5206), .A2(n4465), .ZN(n6854) );
  OAI21_X1 U5246 ( .B1(n6853), .B2(n3874), .A(n6852), .ZN(n2872) );
  NAND2_X1 U5247 ( .A1(n5208), .A2(n4464), .ZN(n6852) );
  OAI21_X1 U5248 ( .B1(n6851), .B2(n3875), .A(n6850), .ZN(n2871) );
  NAND2_X1 U5249 ( .A1(n5207), .A2(n4463), .ZN(n6850) );
  OAI21_X1 U5250 ( .B1(n6832), .B2(n5203), .A(n6831), .ZN(n2864) );
  NAND2_X1 U5251 ( .A1(n5208), .A2(n4249), .ZN(n6831) );
  OAI21_X1 U5252 ( .B1(n6894), .B2(n5204), .A(n6893), .ZN(n2882) );
  NAND2_X1 U5253 ( .A1(n5208), .A2(n4482), .ZN(n6893) );
  OAI21_X1 U5254 ( .B1(n7052), .B2(n5205), .A(n7051), .ZN(n2683) );
  NAND2_X1 U5255 ( .A1(n5206), .A2(\dp/b_adder_id_exe_int[2] ), .ZN(n7051) );
  OAI21_X1 U5256 ( .B1(n7061), .B2(n3874), .A(n7059), .ZN(n2685) );
  NAND2_X1 U5257 ( .A1(n5208), .A2(\dp/b_adder_id_exe_int[0] ), .ZN(n7059) );
  OAI21_X1 U5258 ( .B1(n6889), .B2(n3875), .A(n6888), .ZN(n2881) );
  NAND2_X1 U5259 ( .A1(n5207), .A2(n4255), .ZN(n6888) );
  OAI21_X1 U5260 ( .B1(n6788), .B2(n5203), .A(n6787), .ZN(n2856) );
  NAND2_X1 U5261 ( .A1(n5206), .A2(n4241), .ZN(n6787) );
  OAI21_X1 U5262 ( .B1(n7047), .B2(n5204), .A(n7046), .ZN(n2682) );
  NAND2_X1 U5263 ( .A1(n5208), .A2(\dp/b_adder_id_exe_int[3] ), .ZN(n7046) );
  OAI21_X1 U5264 ( .B1(n6857), .B2(n5205), .A(n6856), .ZN(n2874) );
  NAND2_X1 U5265 ( .A1(n5206), .A2(n4466), .ZN(n6856) );
  OAI211_X1 U5266 ( .C1(n7163), .C2(n4205), .A(n7153), .B(n7161), .ZN(n3056)
         );
  NAND2_X1 U5267 ( .A1(n4097), .A2(rt_id[1]), .ZN(n7153) );
  OAI211_X1 U5268 ( .C1(n7163), .C2(n4258), .A(n7155), .B(n7161), .ZN(n3054)
         );
  NAND2_X1 U5269 ( .A1(n4097), .A2(rt_id[3]), .ZN(n7155) );
  OAI211_X1 U5270 ( .C1(n7163), .C2(n4211), .A(n7162), .B(n7161), .ZN(n3048)
         );
  NAND2_X1 U5271 ( .A1(n4097), .A2(rs_id[4]), .ZN(n7162) );
  NAND2_X1 U5272 ( .A1(n4817), .A2(n6898), .ZN(n2716) );
  AND2_X1 U5273 ( .A1(n6897), .A2(n4334), .ZN(n4817) );
  NAND2_X1 U5274 ( .A1(n3897), .A2(n5146), .ZN(n6897) );
  OAI22_X1 U5275 ( .A1(n6689), .A2(n5196), .B1(n4442), .B2(n5199), .ZN(n2824)
         );
  XNOR2_X1 U5276 ( .A(n6688), .B(n6687), .ZN(n6689) );
  NAND2_X1 U5277 ( .A1(n6686), .A2(n6685), .ZN(n6687) );
  INV_X1 U5278 ( .A(n6682), .ZN(n6683) );
  NAND2_X1 U5279 ( .A1(n6950), .A2(n4819), .ZN(n2701) );
  AND2_X1 U5280 ( .A1(n6949), .A2(n4333), .ZN(n4819) );
  AOI211_X1 U5281 ( .C1(n7436), .C2(rt_id[0]), .A(n6980), .B(n6948), .ZN(n7001) );
  NOR2_X1 U5282 ( .A1(n7004), .A2(n4357), .ZN(n6948) );
  NAND2_X1 U5283 ( .A1(n3896), .A2(n4395), .ZN(n6949) );
  NAND2_X1 U5284 ( .A1(n3956), .A2(\dp/id_exe_regs/b_mult_reg/q[17] ), .ZN(
        n6950) );
  OAI21_X1 U5285 ( .B1(n3935), .B2(n4546), .A(n5547), .ZN(\ctrl_u/n539 ) );
  OAI22_X1 U5286 ( .A1(n6628), .A2(n5196), .B1(n4380), .B2(n5199), .ZN(n2830)
         );
  OAI211_X1 U5287 ( .C1(n6976), .C2(n4582), .A(n6929), .B(n6974), .ZN(n2654)
         );
  NAND2_X1 U5288 ( .A1(n3881), .A2(\dp/ids/rp2[31] ), .ZN(n6929) );
  OAI211_X1 U5289 ( .C1(n6976), .C2(n4293), .A(n6968), .B(n6974), .ZN(n2656)
         );
  NAND2_X1 U5290 ( .A1(n3880), .A2(\dp/ids/rp2[29] ), .ZN(n6968) );
  OAI211_X1 U5291 ( .C1(n6976), .C2(n4291), .A(n6975), .B(n6974), .ZN(n2659)
         );
  NAND2_X1 U5292 ( .A1(n3880), .A2(\dp/ids/rp2[26] ), .ZN(n6975) );
  AOI22_X1 U5293 ( .A1(n5621), .A2(\ctrl_u/next_exe[16] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[16] ), .ZN(\ctrl_u/n445 ) );
  AOI22_X1 U5294 ( .A1(n5621), .A2(\ctrl_u/next_exe[10] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[10] ), .ZN(\ctrl_u/n451 ) );
  AOI22_X1 U5295 ( .A1(n5621), .A2(\ctrl_u/next_exe[12] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[12] ), .ZN(\ctrl_u/n449 ) );
  AOI22_X1 U5296 ( .A1(n5621), .A2(\ctrl_u/next_exe[7] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[7] ), .ZN(\ctrl_u/n454 ) );
  AOI22_X1 U5297 ( .A1(n5621), .A2(\ctrl_u/next_exe[9] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[9] ), .ZN(\ctrl_u/n452 ) );
  AOI22_X1 U5298 ( .A1(n5621), .A2(\ctrl_u/next_exe[14] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[14] ), .ZN(\ctrl_u/n447 ) );
  AOI22_X1 U5299 ( .A1(n5621), .A2(\ctrl_u/next_exe[13] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[13] ), .ZN(\ctrl_u/n448 ) );
  AOI22_X1 U5300 ( .A1(n5621), .A2(\ctrl_u/next_exe[11] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[11] ), .ZN(\ctrl_u/n450 ) );
  AOI22_X1 U5301 ( .A1(n5621), .A2(\ctrl_u/next_exe[8] ), .B1(n5622), .B2(
        \ctrl_u/curr_exe[8] ), .ZN(\ctrl_u/n453 ) );
  OAI22_X1 U5302 ( .A1(n5224), .A2(n4120), .B1(n4362), .B2(n4865), .ZN(n262)
         );
  OAI22_X1 U5303 ( .A1(n5224), .A2(n4501), .B1(n4168), .B2(n4865), .ZN(n252)
         );
  OAI22_X1 U5304 ( .A1(n5224), .A2(n4100), .B1(n4447), .B2(n4865), .ZN(n254)
         );
  OAI22_X1 U5305 ( .A1(n5224), .A2(n4121), .B1(n4372), .B2(n4865), .ZN(n260)
         );
  OAI22_X1 U5306 ( .A1(n5225), .A2(n4118), .B1(n4364), .B2(n4865), .ZN(n264)
         );
  OAI22_X1 U5307 ( .A1(n5225), .A2(\intadd_2/A[0] ), .B1(n4446), .B2(n4865), 
        .ZN(n253) );
  OAI22_X1 U5308 ( .A1(n5225), .A2(\intadd_2/A[2] ), .B1(n4381), .B2(n4865), 
        .ZN(n255) );
  OAI22_X1 U5309 ( .A1(n5225), .A2(n4098), .B1(n4374), .B2(n4865), .ZN(n258)
         );
  OAI22_X1 U5310 ( .A1(n5225), .A2(n4119), .B1(n4363), .B2(n4865), .ZN(n263)
         );
  OAI22_X1 U5311 ( .A1(n5225), .A2(\intadd_2/A[8] ), .B1(n4361), .B2(n4865), 
        .ZN(n261) );
  OAI211_X1 U5312 ( .C1(\intadd_2/SUM[19] ), .C2(n3937), .A(n6399), .B(n6398), 
        .ZN(n2537) );
  AOI22_X1 U5313 ( .A1(n3883), .A2(n6423), .B1(n3928), .B2(
        \dp/pc_plus4_out_if_int[20] ), .ZN(n6398) );
  XNOR2_X1 U5314 ( .A(n4849), .B(n4848), .ZN(\intadd_2/SUM[19] ) );
  XNOR2_X1 U5315 ( .A(n4103), .B(\dp/imm_id_exe_int[22] ), .ZN(n4848) );
  AOI21_X1 U5316 ( .B1(n4032), .B2(n4941), .A(n4826), .ZN(n4849) );
  INV_X1 U5317 ( .A(n4828), .ZN(n4826) );
  NAND2_X1 U5318 ( .A1(n4818), .A2(n6913), .ZN(n2700) );
  NAND2_X1 U5319 ( .A1(n3947), .A2(\dp/id_exe_regs/b_mult_reg/q[18] ), .ZN(
        n6913) );
  AND2_X1 U5320 ( .A1(n6912), .A2(n4332), .ZN(n4818) );
  AOI211_X1 U5321 ( .C1(n7436), .C2(rt_id[1]), .A(n6980), .B(n6911), .ZN(n6996) );
  NOR2_X1 U5322 ( .A1(n6999), .A2(n4357), .ZN(n6911) );
  NAND2_X1 U5323 ( .A1(n3898), .A2(n4394), .ZN(n6912) );
  AOI21_X1 U5324 ( .B1(\dp/ids/rp2[25] ), .B2(b_selector_id), .A(n6920), .ZN(
        n6979) );
  AOI21_X1 U5325 ( .B1(n6919), .B2(n7146), .A(b_selector_id), .ZN(n6920) );
  INV_X1 U5326 ( .A(n6921), .ZN(n6919) );
  OAI211_X1 U5327 ( .C1(n5224), .C2(n4259), .A(n7156), .B(n7161), .ZN(n3053)
         );
  NAND2_X1 U5328 ( .A1(n4097), .A2(rt_id[4]), .ZN(n7156) );
  OAI211_X1 U5329 ( .C1(n5224), .C2(n4221), .A(n7160), .B(n7161), .ZN(n3049)
         );
  NAND2_X1 U5330 ( .A1(n4097), .A2(rs_id[3]), .ZN(n7160) );
  OAI211_X1 U5331 ( .C1(n5224), .C2(n4257), .A(n7154), .B(n7161), .ZN(n3055)
         );
  NAND2_X1 U5332 ( .A1(n4097), .A2(rt_id[2]), .ZN(n7154) );
  OAI211_X1 U5333 ( .C1(n6976), .C2(n4292), .A(n6964), .B(n6974), .ZN(n2655)
         );
  NAND2_X1 U5334 ( .A1(n3880), .A2(\dp/ids/rp2[30] ), .ZN(n6964) );
  OAI211_X1 U5335 ( .C1(n6976), .C2(n4294), .A(n6970), .B(n6974), .ZN(n2657)
         );
  NAND2_X1 U5336 ( .A1(n3881), .A2(\dp/ids/rp2[28] ), .ZN(n6970) );
  OAI211_X1 U5337 ( .C1(n6976), .C2(n4295), .A(n6972), .B(n6974), .ZN(n2658)
         );
  NAND2_X1 U5338 ( .A1(n7005), .A2(n6928), .ZN(n6974) );
  NAND2_X1 U5339 ( .A1(n3881), .A2(\dp/ids/rp2[27] ), .ZN(n6972) );
  INV_X1 U5340 ( .A(n4069), .ZN(n6976) );
  AOI22_X1 U5341 ( .A1(alu_comp_sel[0]), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/next_exe[21] ), .ZN(\ctrl_u/n440 ) );
  AOI22_X1 U5342 ( .A1(op_sign_exe), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/next_exe[27] ), .ZN(\ctrl_u/n434 ) );
  AOI22_X1 U5343 ( .A1(\ctrl_u/curr_exe[20] ), .A2(n5622), .B1(n5621), .B2(
        \ctrl_u/next_exe[20] ), .ZN(\ctrl_u/n441 ) );
  INV_X1 U5344 ( .A(n5137), .ZN(n5676) );
  OAI211_X1 U5345 ( .C1(n5224), .C2(n4220), .A(n7158), .B(n7161), .ZN(n3051)
         );
  NAND2_X1 U5346 ( .A1(n4097), .A2(rs_id[1]), .ZN(n7158) );
  OAI211_X1 U5347 ( .C1(n5224), .C2(n4219), .A(n7152), .B(n7161), .ZN(n3057)
         );
  NAND2_X1 U5348 ( .A1(n4097), .A2(rt_id[0]), .ZN(n7152) );
  OAI211_X1 U5349 ( .C1(n5225), .C2(n3866), .A(n7159), .B(n7161), .ZN(n3050)
         );
  NAND2_X1 U5350 ( .A1(n4097), .A2(rs_id[2]), .ZN(n7159) );
  OAI22_X1 U5351 ( .A1(n6628), .A2(n7062), .B1(n4175), .B2(n3938), .ZN(n2798)
         );
  OAI21_X1 U5352 ( .B1(n5125), .B2(n6630), .A(n6629), .ZN(n6626) );
  NOR2_X1 U5353 ( .A1(n6631), .A2(n6633), .ZN(n6627) );
  OAI211_X1 U5354 ( .C1(n7039), .C2(n4375), .A(n7031), .B(n7030), .ZN(n2678)
         );
  NAND2_X1 U5355 ( .A1(n5209), .A2(\dp/b_adder_id_exe_int[7] ), .ZN(n7030) );
  NAND2_X1 U5356 ( .A1(n3881), .A2(\dp/ids/rp2[7] ), .ZN(n7031) );
  OAI211_X1 U5357 ( .C1(n7039), .C2(n4381), .A(n7038), .B(n7037), .ZN(n2680)
         );
  NAND2_X1 U5358 ( .A1(n5209), .A2(\dp/b_adder_id_exe_int[5] ), .ZN(n7037) );
  NAND2_X1 U5359 ( .A1(n3880), .A2(\dp/ids/rp2[5] ), .ZN(n7038) );
  OAI211_X1 U5360 ( .C1(n7039), .C2(n4376), .A(n7034), .B(n7033), .ZN(n2679)
         );
  NAND2_X1 U5361 ( .A1(n5210), .A2(\dp/b_adder_id_exe_int[6] ), .ZN(n7033) );
  NAND2_X1 U5362 ( .A1(n3880), .A2(\dp/ids/rp2[6] ), .ZN(n7034) );
  OAI211_X1 U5363 ( .C1(n5225), .C2(n4222), .A(n7157), .B(n7161), .ZN(n3052)
         );
  INV_X1 U5364 ( .A(n7146), .ZN(n7150) );
  NAND2_X1 U5365 ( .A1(n4097), .A2(rs_id[0]), .ZN(n7157) );
  OAI22_X1 U5366 ( .A1(n6668), .A2(n5196), .B1(n4387), .B2(n5199), .ZN(n2826)
         );
  OAI21_X1 U5367 ( .B1(n3935), .B2(\ctrl_u/n63 ), .A(n5571), .ZN(\ctrl_u/n513 ) );
  NAND2_X1 U5368 ( .A1(n5646), .A2(n5590), .ZN(n5567) );
  OAI21_X1 U5369 ( .B1(n5182), .B2(n5566), .A(n5571), .ZN(\ctrl_u/n553 ) );
  OAI22_X1 U5370 ( .A1(n6566), .A2(n5197), .B1(n4405), .B2(n5199), .ZN(n2838)
         );
  OAI21_X1 U5371 ( .B1(n5182), .B2(\ctrl_u/n65 ), .A(n5571), .ZN(\ctrl_u/n517 ) );
  OAI211_X1 U5372 ( .C1(n7039), .C2(n4364), .A(n7010), .B(n7009), .ZN(n2671)
         );
  NAND2_X1 U5373 ( .A1(n5210), .A2(\dp/b_adder_id_exe_int[14] ), .ZN(n7009) );
  NAND2_X1 U5374 ( .A1(n3881), .A2(\dp/ids/rp2[14] ), .ZN(n7010) );
  AOI22_X1 U5375 ( .A1(n5134), .A2(\dp/imm_id_int[6] ), .B1(n5180), .B2(
        instr_if[6]), .ZN(n1636) );
  AOI22_X1 U5376 ( .A1(n5134), .A2(\ctrl_u/curr_pt_id ), .B1(n5180), .B2(
        predicted_taken), .ZN(\ctrl_u/n167 ) );
  OAI22_X1 U5377 ( .A1(n6476), .A2(n5197), .B1(n4403), .B2(n5199), .ZN(n2850)
         );
  NOR2_X1 U5378 ( .A1(n6474), .A2(n6479), .ZN(n6475) );
  INV_X1 U5379 ( .A(n6480), .ZN(n6474) );
  OAI22_X1 U5380 ( .A1(n6495), .A2(n5196), .B1(n4453), .B2(n5199), .ZN(n2847)
         );
  INV_X1 U5381 ( .A(n6492), .ZN(n6494) );
  OAI21_X1 U5382 ( .B1(n6701), .B2(n4329), .A(n4913), .ZN(n4912) );
  AOI21_X1 U5383 ( .B1(n6490), .B2(n6491), .A(n6489), .ZN(n4913) );
  INV_X1 U5384 ( .A(n6486), .ZN(n6487) );
  AOI22_X1 U5385 ( .A1(n5133), .A2(\dp/imm_id_int[14] ), .B1(n5179), .B2(
        instr_if[14]), .ZN(n1628) );
  AOI22_X1 U5386 ( .A1(n5133), .A2(\dp/imm_id_int[13] ), .B1(n3978), .B2(
        instr_if[13]), .ZN(n1629) );
  AOI22_X1 U5387 ( .A1(n5133), .A2(\dp/imm_id_int[15] ), .B1(n5179), .B2(
        instr_if[15]), .ZN(n1627) );
  OAI22_X1 U5388 ( .A1(n6517), .A2(n5196), .B1(n4474), .B2(n5199), .ZN(n2844)
         );
  OAI211_X1 U5389 ( .C1(n4368), .C2(n7039), .A(n7007), .B(n7006), .ZN(n2670)
         );
  NAND2_X1 U5390 ( .A1(n5209), .A2(\dp/b_adder_id_exe_int[15] ), .ZN(n7006) );
  NAND2_X1 U5391 ( .A1(n3880), .A2(\dp/ids/rp2[15] ), .ZN(n7007) );
  OR2_X1 U5392 ( .A1(n5443), .A2(n5619), .ZN(\ctrl_u/n536 ) );
  OAI21_X1 U5393 ( .B1(n5440), .B2(n5439), .A(n5502), .ZN(n5441) );
  OAI211_X1 U5394 ( .C1(n5494), .C2(n5560), .A(n5650), .B(n5514), .ZN(n5439)
         );
  OAI21_X1 U5395 ( .B1(n3934), .B2(n4545), .A(n3857), .ZN(\ctrl_u/n538 ) );
  OAI211_X1 U5396 ( .C1(n3935), .C2(n4579), .A(n5547), .B(n5488), .ZN(
        \ctrl_u/n505 ) );
  OAI21_X1 U5397 ( .B1(n5182), .B2(\ctrl_u/n67 ), .A(n5570), .ZN(\ctrl_u/n519 ) );
  OAI22_X1 U5398 ( .A1(n5219), .A2(n373), .B1(n3891), .B2(n4207), .ZN(n2995)
         );
  OAI22_X1 U5399 ( .A1(n5218), .A2(n365), .B1(n3892), .B2(n4210), .ZN(n3003)
         );
  OAI22_X1 U5400 ( .A1(n5222), .A2(n383), .B1(n3889), .B2(n4137), .ZN(n2985)
         );
  OAI22_X1 U5401 ( .A1(n5223), .A2(n367), .B1(n3893), .B2(n4217), .ZN(n3001)
         );
  OAI22_X1 U5402 ( .A1(n5222), .A2(n389), .B1(n3893), .B2(n4483), .ZN(n2979)
         );
  OAI22_X1 U5403 ( .A1(n5218), .A2(n381), .B1(n3891), .B2(\intadd_2/B[20] ), 
        .ZN(n2987) );
  OAI22_X1 U5404 ( .A1(n5223), .A2(n374), .B1(n3893), .B2(n4102), .ZN(n2994)
         );
  OAI22_X1 U5405 ( .A1(n5221), .A2(n375), .B1(n3893), .B2(\intadd_2/B[14] ), 
        .ZN(n2993) );
  OAI21_X1 U5406 ( .B1(n5182), .B2(\ctrl_u/n68 ), .A(n3857), .ZN(\ctrl_u/n520 ) );
  OAI22_X1 U5407 ( .A1(n5563), .A2(n5559), .B1(n3935), .B2(n4541), .ZN(
        \ctrl_u/n546 ) );
  INV_X1 U5408 ( .A(n5558), .ZN(n5559) );
  OAI211_X1 U5409 ( .C1(n7039), .C2(n4361), .A(n7019), .B(n7018), .ZN(n2674)
         );
  NAND2_X1 U5410 ( .A1(n5207), .A2(\dp/b_adder_id_exe_int[11] ), .ZN(n7018) );
  NAND2_X1 U5411 ( .A1(n3881), .A2(\dp/ids/rp2[11] ), .ZN(n7019) );
  OAI211_X1 U5412 ( .C1(n7039), .C2(n4373), .A(n7025), .B(n7024), .ZN(n2676)
         );
  NAND2_X1 U5413 ( .A1(n5207), .A2(\dp/b_adder_id_exe_int[9] ), .ZN(n7024) );
  NAND2_X1 U5414 ( .A1(n3880), .A2(\dp/ids/rp2[9] ), .ZN(n7025) );
  OAI211_X1 U5415 ( .C1(n7039), .C2(n4363), .A(n7013), .B(n7012), .ZN(n2672)
         );
  NAND2_X1 U5416 ( .A1(n5208), .A2(\dp/b_adder_id_exe_int[13] ), .ZN(n7012) );
  NAND2_X1 U5417 ( .A1(n3881), .A2(\dp/ids/rp2[13] ), .ZN(n7013) );
  OAI211_X1 U5418 ( .C1(n7039), .C2(n4374), .A(n7028), .B(n7027), .ZN(n2677)
         );
  NAND2_X1 U5419 ( .A1(n5208), .A2(\dp/b_adder_id_exe_int[8] ), .ZN(n7027) );
  NAND2_X1 U5420 ( .A1(n3880), .A2(\dp/ids/rp2[8] ), .ZN(n7028) );
  OAI211_X1 U5421 ( .C1(n7039), .C2(n4372), .A(n7022), .B(n7021), .ZN(n2675)
         );
  NAND2_X1 U5422 ( .A1(n5208), .A2(\dp/b_adder_id_exe_int[10] ), .ZN(n7021) );
  NAND2_X1 U5423 ( .A1(n3881), .A2(\dp/ids/rp2[10] ), .ZN(n7022) );
  OAI211_X1 U5424 ( .C1(n7039), .C2(n4362), .A(n7016), .B(n7015), .ZN(n2673)
         );
  NAND2_X1 U5425 ( .A1(n5206), .A2(\dp/b_adder_id_exe_int[12] ), .ZN(n7015) );
  NAND2_X1 U5426 ( .A1(n3880), .A2(\dp/ids/rp2[12] ), .ZN(n7016) );
  AOI21_X1 U5427 ( .B1(rp2_out_sel_id[0]), .B2(n3941), .A(n5489), .ZN(
        \ctrl_u/n181 ) );
  AOI21_X1 U5428 ( .B1(rp2_out_sel_id[1]), .B2(n3941), .A(n5489), .ZN(
        \ctrl_u/n179 ) );
  NOR2_X1 U5429 ( .A1(n5627), .A2(n5430), .ZN(n5481) );
  INV_X1 U5430 ( .A(n6947), .ZN(n4675) );
  AOI22_X1 U5431 ( .A1(n3896), .A2(\dp/id_exe_regs/b_mult_reg/q[25] ), .B1(
        n3956), .B2(\dp/id_exe_regs/b_mult_reg/q[27] ), .ZN(n6959) );
  NAND2_X1 U5432 ( .A1(n5214), .A2(\dp/ids/rp2[26] ), .ZN(n6960) );
  OAI22_X1 U5433 ( .A1(n6668), .A2(n7062), .B1(n4187), .B2(n3938), .ZN(n2794)
         );
  OAI21_X1 U5434 ( .B1(n6701), .B2(n6670), .A(n6669), .ZN(n6666) );
  NOR2_X1 U5435 ( .A1(n6671), .A2(n6673), .ZN(n6667) );
  OAI22_X1 U5436 ( .A1(n6559), .A2(n5196), .B1(n4475), .B2(n5199), .ZN(n2839)
         );
  OAI22_X1 U5437 ( .A1(n6517), .A2(n7062), .B1(n4183), .B2(n3938), .ZN(n2812)
         );
  OAI21_X1 U5438 ( .B1(n6701), .B2(n6521), .A(n6520), .ZN(n6515) );
  NOR2_X1 U5439 ( .A1(n6522), .A2(n6524), .ZN(n6516) );
  OAI22_X1 U5440 ( .A1(n6566), .A2(n7062), .B1(n4173), .B2(n3938), .ZN(n2806)
         );
  OAI21_X1 U5441 ( .B1(n6701), .B2(n6578), .A(n6581), .ZN(n6564) );
  NOR2_X1 U5442 ( .A1(n6567), .A2(n6569), .ZN(n6565) );
  OAI22_X1 U5443 ( .A1(n6710), .A2(n5198), .B1(n4452), .B2(n5199), .ZN(n2821)
         );
  AOI22_X1 U5444 ( .A1(n5134), .A2(\dp/imm_id_int[1] ), .B1(n5179), .B2(
        instr_if[1]), .ZN(n1641) );
  AOI22_X1 U5445 ( .A1(n5134), .A2(\dp/imm_id_int[3] ), .B1(n5179), .B2(
        instr_if[3]), .ZN(n1639) );
  AOI22_X1 U5446 ( .A1(n5134), .A2(\dp/imm_id_int[2] ), .B1(n5179), .B2(
        instr_if[2]), .ZN(n1640) );
  AOI22_X1 U5447 ( .A1(n5133), .A2(\dp/imm_id_int[9] ), .B1(n5179), .B2(
        instr_if[9]), .ZN(n1633) );
  AOI22_X1 U5448 ( .A1(n5133), .A2(\dp/imm_id_int[10] ), .B1(n5179), .B2(
        instr_if[10]), .ZN(n1632) );
  AOI22_X1 U5449 ( .A1(n5133), .A2(\dp/imm_id_int[11] ), .B1(n5179), .B2(
        instr_if[11]), .ZN(n1631) );
  OAI211_X1 U5450 ( .C1(n4359), .C2(n7170), .A(n7169), .B(n7168), .ZN(n3063)
         );
  AOI22_X1 U5451 ( .A1(n7167), .A2(\dp/imm_id_int[15] ), .B1(n7166), .B2(
        rd_idexe[4]), .ZN(n7169) );
  INV_X1 U5452 ( .A(n7165), .ZN(n7167) );
  INV_X1 U5453 ( .A(n7164), .ZN(n7170) );
  OAI22_X1 U5454 ( .A1(n6559), .A2(n7062), .B1(n4185), .B2(n3942), .ZN(n2807)
         );
  XNOR2_X1 U5455 ( .A(n6558), .B(n6557), .ZN(n6559) );
  NOR2_X1 U5456 ( .A1(n6556), .A2(n6555), .ZN(n6557) );
  INV_X1 U5457 ( .A(n6554), .ZN(n6556) );
  INV_X1 U5458 ( .A(n6547), .ZN(n6552) );
  OAI22_X1 U5459 ( .A1(n6710), .A2(n7062), .B1(n4179), .B2(n3942), .ZN(n2789)
         );
  XNOR2_X1 U5460 ( .A(n6709), .B(n6708), .ZN(n6710) );
  NOR2_X1 U5461 ( .A1(n6707), .A2(n6706), .ZN(n6708) );
  OAI22_X1 U5462 ( .A1(n6577), .A2(n7062), .B1(n4174), .B2(n3942), .ZN(n2805)
         );
  OAI22_X1 U5463 ( .A1(n6546), .A2(n7062), .B1(n4184), .B2(n3938), .ZN(n2808)
         );
  OAI21_X1 U5464 ( .B1(n6681), .B2(n5196), .A(n4809), .ZN(n2825) );
  NAND2_X1 U5465 ( .A1(n7098), .A2(\dp/a_neg_mult_id_exe_int[57] ), .ZN(n4809)
         );
  OAI22_X1 U5466 ( .A1(n6698), .A2(n5197), .B1(n4451), .B2(n4808), .ZN(n2822)
         );
  OAI22_X1 U5467 ( .A1(n5196), .A2(n6546), .B1(n4471), .B2(n4808), .ZN(n2840)
         );
  AOI21_X1 U5468 ( .B1(n6563), .B2(n6543), .A(n6542), .ZN(n6547) );
  NAND2_X1 U5469 ( .A1(n6560), .A2(n6543), .ZN(n6548) );
  INV_X1 U5470 ( .A(n6541), .ZN(n6543) );
  NOR2_X1 U5471 ( .A1(n6549), .A2(n6551), .ZN(n6545) );
  INV_X1 U5472 ( .A(n6553), .ZN(n6549) );
  OAI22_X1 U5473 ( .A1(n5218), .A2(n360), .B1(n3889), .B2(
        btb_cache_rw_address[0]), .ZN(n3008) );
  OAI22_X1 U5474 ( .A1(n5221), .A2(n382), .B1(n3890), .B2(n4356), .ZN(n2986)
         );
  OAI22_X1 U5475 ( .A1(n5219), .A2(n380), .B1(n3890), .B2(n4103), .ZN(n2988)
         );
  OAI22_X1 U5476 ( .A1(n5219), .A2(n379), .B1(n3891), .B2(n4101), .ZN(n2989)
         );
  OAI22_X1 U5477 ( .A1(n5218), .A2(n378), .B1(n3891), .B2(n4114), .ZN(n2990)
         );
  OAI22_X1 U5478 ( .A1(n5223), .A2(n377), .B1(n3892), .B2(n4110), .ZN(n2991)
         );
  OAI22_X1 U5479 ( .A1(n5222), .A2(n376), .B1(n3892), .B2(n4113), .ZN(n2992)
         );
  OAI22_X1 U5480 ( .A1(n5221), .A2(n388), .B1(n3891), .B2(n4519), .ZN(n2980)
         );
  OAI22_X1 U5481 ( .A1(n5222), .A2(n371), .B1(n3892), .B2(n4226), .ZN(n2997)
         );
  OAI22_X1 U5482 ( .A1(n5220), .A2(n387), .B1(n3893), .B2(n4536), .ZN(n2981)
         );
  OAI22_X1 U5483 ( .A1(n5220), .A2(n386), .B1(n3893), .B2(n4148), .ZN(n2982)
         );
  OAI22_X1 U5484 ( .A1(n5222), .A2(n361), .B1(n3892), .B2(n4213), .ZN(n3007)
         );
  OAI22_X1 U5485 ( .A1(n5220), .A2(n385), .B1(n3890), .B2(n4520), .ZN(n2983)
         );
  OAI22_X1 U5486 ( .A1(n5223), .A2(n384), .B1(n3890), .B2(n4147), .ZN(n2984)
         );
  OAI22_X1 U5487 ( .A1(n5220), .A2(n364), .B1(n3889), .B2(n4215), .ZN(n3004)
         );
  OAI22_X1 U5488 ( .A1(n5219), .A2(n363), .B1(n3893), .B2(n4209), .ZN(n3005)
         );
  OAI22_X1 U5489 ( .A1(n5219), .A2(n362), .B1(n3890), .B2(n4214), .ZN(n3006)
         );
  OAI22_X1 U5490 ( .A1(n5221), .A2(n369), .B1(n3889), .B2(n4218), .ZN(n2999)
         );
  OAI22_X1 U5491 ( .A1(n5221), .A2(n370), .B1(n3889), .B2(n4234), .ZN(n2998)
         );
  OAI22_X1 U5492 ( .A1(n5220), .A2(n368), .B1(n3893), .B2(n4233), .ZN(n3000)
         );
  OAI22_X1 U5493 ( .A1(n5223), .A2(n372), .B1(n3889), .B2(n4235), .ZN(n2996)
         );
  OAI22_X1 U5494 ( .A1(n5218), .A2(n366), .B1(n3890), .B2(n4216), .ZN(n3002)
         );
  NOR2_X1 U5495 ( .A1(n6716), .A2(n6715), .ZN(n6717) );
  INV_X1 U5496 ( .A(n6711), .ZN(n6713) );
  NOR2_X1 U5497 ( .A1(n6488), .A2(n6489), .ZN(n6483) );
  INV_X1 U5498 ( .A(n6491), .ZN(n6488) );
  NOR2_X1 U5499 ( .A1(n6582), .A2(n6587), .ZN(n6583) );
  INV_X1 U5500 ( .A(n6589), .ZN(n6582) );
  OAI21_X1 U5501 ( .B1(n6581), .B2(n6580), .A(n6579), .ZN(n6588) );
  NOR2_X1 U5502 ( .A1(n6578), .A2(n6580), .ZN(n6586) );
  OAI211_X1 U5503 ( .C1(\intadd_2/SUM[18] ), .C2(n3937), .A(n6397), .B(n6396), 
        .ZN(n2538) );
  AOI22_X1 U5504 ( .A1(n3883), .A2(n6425), .B1(n3936), .B2(
        \dp/pc_plus4_out_if_int[19] ), .ZN(n6396) );
  OAI21_X1 U5505 ( .B1(n6018), .B2(n6027), .A(n6017), .ZN(n6425) );
  AOI21_X1 U5506 ( .B1(\dp/exs/alu_unit/shifter_out[21] ), .B2(n7083), .A(
        n6016), .ZN(n6017) );
  OAI21_X1 U5507 ( .B1(\intadd_1/SUM[20] ), .B2(n7066), .A(n6015), .ZN(n6016)
         );
  NAND2_X1 U5508 ( .A1(n6012), .A2(n3952), .ZN(n6013) );
  NAND2_X1 U5509 ( .A1(n4862), .A2(n4902), .ZN(n6022) );
  NAND2_X1 U5510 ( .A1(n5988), .A2(n4904), .ZN(n4862) );
  INV_X1 U5511 ( .A(n6395), .ZN(n6397) );
  XNOR2_X1 U5512 ( .A(n4032), .B(n4942), .ZN(\intadd_2/SUM[18] ) );
  XNOR2_X1 U5513 ( .A(n4101), .B(n4222), .ZN(n4942) );
  OAI211_X1 U5514 ( .C1(n3873), .C2(n4215), .A(n6351), .B(n6350), .ZN(n2553)
         );
  AOI22_X1 U5515 ( .A1(n3894), .A2(\dp/ifs/pc_btb[4] ), .B1(n5193), .B2(
        btb_cache_read_address[4]), .ZN(n6350) );
  AOI211_X1 U5516 ( .C1(n3936), .C2(\dp/pc_plus4_out_if_int[4] ), .A(n6349), 
        .B(n6348), .ZN(n6351) );
  AND2_X1 U5517 ( .A1(n3884), .A2(n4884), .ZN(n6348) );
  AOI21_X1 U5518 ( .B1(\dp/exs/alu_unit/shifter_out[6] ), .B2(n3954), .A(n5880), .ZN(n6457) );
  OAI211_X1 U5519 ( .C1(\intadd_1/SUM[5] ), .C2(n7066), .A(n5879), .B(n5878), 
        .ZN(n5880) );
  NAND2_X1 U5520 ( .A1(n5877), .A2(n7076), .ZN(n5878) );
  XNOR2_X1 U5521 ( .A(n5876), .B(n5875), .ZN(n5877) );
  AOI21_X1 U5522 ( .B1(n5873), .B2(n5872), .A(n5871), .ZN(n5876) );
  INV_X1 U5523 ( .A(n5872), .ZN(n5869) );
  INV_X1 U5524 ( .A(n5870), .ZN(n5873) );
  NAND2_X1 U5525 ( .A1(n5865), .A2(n3952), .ZN(n5866) );
  NOR2_X1 U5526 ( .A1(n3879), .A2(\intadd_2/SUM[3] ), .ZN(n6349) );
  XNOR2_X1 U5527 ( .A(n5075), .B(n5074), .ZN(\intadd_2/SUM[3] ) );
  XNOR2_X1 U5528 ( .A(n4215), .B(n4099), .ZN(n5074) );
  OAI211_X1 U5529 ( .C1(n3873), .C2(n4210), .A(n6355), .B(n6354), .ZN(n2552)
         );
  AOI22_X1 U5530 ( .A1(n3931), .A2(\dp/ifs/pc_btb[5] ), .B1(n5193), .B2(
        btb_cache_read_address[5]), .ZN(n6354) );
  AOI211_X1 U5531 ( .C1(n3928), .C2(\dp/pc_plus4_out_if_int[5] ), .A(n6353), 
        .B(n6352), .ZN(n6355) );
  AND2_X1 U5532 ( .A1(n3884), .A2(n4885), .ZN(n6352) );
  OAI211_X1 U5533 ( .C1(\intadd_1/SUM[6] ), .C2(n7066), .A(n5891), .B(n5890), 
        .ZN(n5892) );
  NAND2_X1 U5534 ( .A1(n5889), .A2(n7076), .ZN(n5890) );
  XNOR2_X1 U5535 ( .A(n5886), .B(n5885), .ZN(n5887) );
  NAND2_X1 U5536 ( .A1(n4042), .A2(n3952), .ZN(n5883) );
  NOR2_X1 U5537 ( .A1(n3879), .A2(\intadd_2/SUM[4] ), .ZN(n6353) );
  OAI211_X1 U5538 ( .C1(n3873), .C2(n4213), .A(n6339), .B(n6338), .ZN(n2556)
         );
  AOI22_X1 U5539 ( .A1(n3894), .A2(\dp/ifs/pc_btb[1] ), .B1(n5193), .B2(
        btb_cache_read_address[1]), .ZN(n6338) );
  AOI211_X1 U5540 ( .C1(n3936), .C2(\dp/pc_plus4_out_if_int[1] ), .A(n6337), 
        .B(n6336), .ZN(n6339) );
  AND2_X1 U5541 ( .A1(n3884), .A2(n4881), .ZN(n6336) );
  OAI211_X1 U5542 ( .C1(\intadd_1/SUM[2] ), .C2(n7066), .A(n5834), .B(n5833), 
        .ZN(n5835) );
  NAND2_X1 U5543 ( .A1(n5832), .A2(n7076), .ZN(n5833) );
  XNOR2_X1 U5544 ( .A(n5831), .B(n5842), .ZN(n5832) );
  XNOR2_X1 U5545 ( .A(n5841), .B(n5840), .ZN(n5831) );
  NAND2_X1 U5546 ( .A1(n5828), .A2(n3952), .ZN(n5829) );
  NOR2_X1 U5547 ( .A1(n3879), .A2(\intadd_2/SUM[0] ), .ZN(n6337) );
  XNOR2_X1 U5548 ( .A(n4213), .B(n5094), .ZN(\intadd_2/SUM[0] ) );
  XNOR2_X1 U5549 ( .A(n5095), .B(\intadd_2/A[0] ), .ZN(n5094) );
  OAI211_X1 U5550 ( .C1(n3873), .C2(n4216), .A(n6359), .B(n6358), .ZN(n2551)
         );
  AOI22_X1 U5551 ( .A1(n3895), .A2(\dp/ifs/pc_btb[6] ), .B1(n5193), .B2(
        btb_cache_read_address[6]), .ZN(n6358) );
  AOI211_X1 U5552 ( .C1(n3928), .C2(\dp/pc_plus4_out_if_int[6] ), .A(n6357), 
        .B(n6356), .ZN(n6359) );
  AND2_X1 U5553 ( .A1(n3884), .A2(n4886), .ZN(n6356) );
  AOI21_X1 U5554 ( .B1(\dp/exs/alu_unit/shifter_out[8] ), .B2(n3954), .A(n5904), .ZN(n6451) );
  OAI211_X1 U5555 ( .C1(\intadd_1/SUM[7] ), .C2(n7066), .A(n5903), .B(n5902), 
        .ZN(n5904) );
  NAND2_X1 U5556 ( .A1(n5901), .A2(n7076), .ZN(n5902) );
  NAND2_X1 U5557 ( .A1(n5112), .A2(n3952), .ZN(n5895) );
  INV_X1 U5558 ( .A(n5894), .ZN(n5112) );
  NOR2_X1 U5559 ( .A1(n3879), .A2(\intadd_2/SUM[5] ), .ZN(n6357) );
  XNOR2_X1 U5560 ( .A(n5022), .B(n5021), .ZN(\intadd_2/SUM[5] ) );
  XNOR2_X1 U5561 ( .A(n4216), .B(n4098), .ZN(n5021) );
  NAND2_X1 U5562 ( .A1(n5000), .A2(n5039), .ZN(n5022) );
  NAND2_X1 U5563 ( .A1(n5075), .A2(n5040), .ZN(n5000) );
  OAI211_X1 U5564 ( .C1(n3873), .C2(n4217), .A(n6363), .B(n6362), .ZN(n2550)
         );
  AOI22_X1 U5565 ( .A1(n3895), .A2(\dp/ifs/pc_btb[7] ), .B1(n5193), .B2(
        btb_cache_read_address[7]), .ZN(n6362) );
  AOI211_X1 U5566 ( .C1(n3928), .C2(\dp/pc_plus4_out_if_int[7] ), .A(n6361), 
        .B(n6360), .ZN(n6363) );
  AND2_X1 U5567 ( .A1(n3884), .A2(n4887), .ZN(n6360) );
  AOI21_X1 U5568 ( .B1(\dp/exs/alu_unit/shifter_out[9] ), .B2(n3954), .A(n5915), .ZN(n6449) );
  OAI211_X1 U5569 ( .C1(\intadd_1/SUM[8] ), .C2(n7066), .A(n5914), .B(n5913), 
        .ZN(n5915) );
  NAND2_X1 U5570 ( .A1(n5912), .A2(n7076), .ZN(n5913) );
  XNOR2_X1 U5571 ( .A(n5909), .B(n5908), .ZN(n5910) );
  NAND2_X1 U5572 ( .A1(n5115), .A2(n3952), .ZN(n5906) );
  INV_X1 U5573 ( .A(n4672), .ZN(n5115) );
  BUF_X1 U5574 ( .A(n5144), .Z(n4672) );
  NOR2_X1 U5575 ( .A1(n3879), .A2(\intadd_2/SUM[6] ), .ZN(n6361) );
  OAI211_X1 U5576 ( .C1(n3873), .C2(n4214), .A(n6343), .B(n6342), .ZN(n2555)
         );
  AOI22_X1 U5577 ( .A1(n3895), .A2(\dp/ifs/pc_btb[2] ), .B1(n5193), .B2(
        btb_cache_read_address[2]), .ZN(n6342) );
  AOI211_X1 U5578 ( .C1(n3936), .C2(\dp/pc_plus4_out_if_int[2] ), .A(n6341), 
        .B(n6340), .ZN(n6343) );
  AND2_X1 U5579 ( .A1(n3884), .A2(n4882), .ZN(n6340) );
  AOI21_X1 U5580 ( .B1(\dp/exs/alu_unit/shifter_out[4] ), .B2(n7083), .A(n5849), .ZN(n6462) );
  OAI211_X1 U5581 ( .C1(\intadd_1/SUM[3] ), .C2(n7066), .A(n5848), .B(n5847), 
        .ZN(n5849) );
  NAND2_X1 U5582 ( .A1(n5846), .A2(n7076), .ZN(n5847) );
  XNOR2_X1 U5583 ( .A(n5856), .B(n5845), .ZN(n5846) );
  NAND2_X1 U5584 ( .A1(n5114), .A2(n3940), .ZN(n5838) );
  INV_X1 U5585 ( .A(\intadd_1/B[3] ), .ZN(n5114) );
  NOR2_X1 U5586 ( .A1(n3879), .A2(\intadd_2/SUM[1] ), .ZN(n6341) );
  XNOR2_X1 U5587 ( .A(n5084), .B(n5083), .ZN(\intadd_2/SUM[1] ) );
  XNOR2_X1 U5588 ( .A(n4214), .B(n4100), .ZN(n5083) );
  OAI211_X1 U5589 ( .C1(n3873), .C2(n4233), .A(n6367), .B(n6366), .ZN(n2549)
         );
  AOI22_X1 U5590 ( .A1(n3931), .A2(\dp/ifs/pc_btb[8] ), .B1(n7108), .B2(
        btb_cache_read_address[8]), .ZN(n6366) );
  AOI211_X1 U5591 ( .C1(n3936), .C2(\dp/pc_plus4_out_if_int[8] ), .A(n6365), 
        .B(n6364), .ZN(n6367) );
  AND2_X1 U5592 ( .A1(n3884), .A2(n4888), .ZN(n6364) );
  NOR2_X1 U5593 ( .A1(n3879), .A2(\intadd_2/SUM[7] ), .ZN(n6365) );
  OAI211_X1 U5594 ( .C1(n3873), .C2(n4218), .A(n6371), .B(n6370), .ZN(n2548)
         );
  AOI22_X1 U5595 ( .A1(n3894), .A2(\dp/ifs/pc_btb[9] ), .B1(n5193), .B2(
        btb_cache_read_address[9]), .ZN(n6370) );
  AOI211_X1 U5596 ( .C1(n3936), .C2(\dp/pc_plus4_out_if_int[9] ), .A(n6369), 
        .B(n6368), .ZN(n6371) );
  AND2_X1 U5597 ( .A1(n3884), .A2(n4889), .ZN(n6368) );
  NOR2_X1 U5598 ( .A1(n3879), .A2(\intadd_2/SUM[8] ), .ZN(n6369) );
  NOR2_X1 U5599 ( .A1(n6535), .A2(n6537), .ZN(n6529) );
  OAI211_X1 U5600 ( .C1(n3873), .C2(n4209), .A(n6347), .B(n6346), .ZN(n2554)
         );
  AOI22_X1 U5601 ( .A1(n3894), .A2(\dp/ifs/pc_btb[3] ), .B1(n7108), .B2(
        btb_cache_read_address[3]), .ZN(n6346) );
  AOI211_X1 U5602 ( .C1(n3928), .C2(\dp/pc_plus4_out_if_int[3] ), .A(n6345), 
        .B(n6344), .ZN(n6347) );
  AND2_X1 U5603 ( .A1(n3884), .A2(n4883), .ZN(n6344) );
  OAI211_X1 U5604 ( .C1(n4995), .C2(n7066), .A(n5862), .B(n5861), .ZN(n5863)
         );
  NAND2_X1 U5605 ( .A1(n5860), .A2(n7076), .ZN(n5861) );
  XNOR2_X1 U5606 ( .A(n5870), .B(n5859), .ZN(n5860) );
  INV_X1 U5607 ( .A(n5856), .ZN(n5858) );
  NAND2_X1 U5608 ( .A1(n5844), .A2(n5843), .ZN(n5856) );
  NAND2_X1 U5609 ( .A1(n5842), .A2(n5841), .ZN(n5843) );
  OAI21_X1 U5610 ( .B1(n5842), .B2(n5841), .A(n5840), .ZN(n5844) );
  NAND2_X1 U5611 ( .A1(n5851), .A2(n3952), .ZN(n5852) );
  NOR2_X1 U5612 ( .A1(n4734), .A2(n5260), .ZN(n5851) );
  NOR2_X1 U5613 ( .A1(n3879), .A2(\intadd_2/SUM[2] ), .ZN(n6345) );
  XNOR2_X1 U5614 ( .A(n5080), .B(n5079), .ZN(\intadd_2/SUM[2] ) );
  XNOR2_X1 U5615 ( .A(n4209), .B(\intadd_2/A[2] ), .ZN(n5079) );
  OAI21_X1 U5616 ( .B1(n5056), .B2(n4129), .A(n5082), .ZN(n5080) );
  INV_X1 U5617 ( .A(n5084), .ZN(n5056) );
  NOR2_X1 U5618 ( .A1(n6608), .A2(n6613), .ZN(n6609) );
  INV_X1 U5619 ( .A(n6615), .ZN(n6608) );
  OAI211_X1 U5620 ( .C1(n3873), .C2(n4102), .A(n6385), .B(n6384), .ZN(n2543)
         );
  AOI22_X1 U5621 ( .A1(n3931), .A2(\dp/ifs/pc_btb[14] ), .B1(n5193), .B2(
        btb_cache_read_address[14]), .ZN(n6384) );
  AOI211_X1 U5622 ( .C1(n3936), .C2(\dp/pc_plus4_out_if_int[14] ), .A(n6383), 
        .B(n6382), .ZN(n6385) );
  AND2_X1 U5623 ( .A1(n3884), .A2(n4891), .ZN(n6382) );
  NOR2_X1 U5624 ( .A1(n3879), .A2(\intadd_2/SUM[13] ), .ZN(n6383) );
  XNOR2_X1 U5625 ( .A(n4949), .B(n4948), .ZN(\intadd_2/SUM[13] ) );
  XNOR2_X1 U5626 ( .A(n4102), .B(\dp/imm_id_exe_int[16] ), .ZN(n4948) );
  AOI21_X1 U5627 ( .B1(\intadd_2/n17 ), .B2(n5002), .A(n4928), .ZN(n4949) );
  INV_X1 U5628 ( .A(n4930), .ZN(n4928) );
  AOI22_X1 U5629 ( .A1(n3897), .A2(\dp/id_exe_regs/b_mult_reg/q[28] ), .B1(
        n3956), .B2(\dp/id_exe_regs/b_mult_reg/q[30] ), .ZN(n6926) );
  NAND2_X1 U5630 ( .A1(n5213), .A2(\dp/ids/rp2[29] ), .ZN(n6927) );
  OAI211_X1 U5631 ( .C1(n3873), .C2(n4207), .A(n6381), .B(n6380), .ZN(n2544)
         );
  AOI22_X1 U5632 ( .A1(n3894), .A2(\dp/ifs/pc_btb[13] ), .B1(n5193), .B2(
        btb_cache_read_address[13]), .ZN(n6380) );
  AOI211_X1 U5633 ( .C1(n3928), .C2(\dp/pc_plus4_out_if_int[13] ), .A(n6379), 
        .B(n6378), .ZN(n6381) );
  AND2_X1 U5634 ( .A1(n3884), .A2(n4890), .ZN(n6378) );
  AOI21_X1 U5635 ( .B1(n7076), .B2(n5951), .A(n5950), .ZN(n6434) );
  NAND2_X1 U5636 ( .A1(\dp/exs/alu_unit/shifter_out[15] ), .A2(n3954), .ZN(
        n5948) );
  NAND2_X1 U5637 ( .A1(n5116), .A2(n3952), .ZN(n5946) );
  OAI21_X1 U5638 ( .B1(n5116), .B2(n3940), .A(n5008), .ZN(n5947) );
  NAND2_X1 U5639 ( .A1(n5116), .A2(n7069), .ZN(n5008) );
  XNOR2_X1 U5640 ( .A(n5943), .B(n5942), .ZN(n5944) );
  NOR2_X1 U5641 ( .A1(n3879), .A2(\intadd_2/SUM[12] ), .ZN(n6379) );
  XNOR2_X1 U5642 ( .A(\intadd_2/n17 ), .B(n5003), .ZN(\intadd_2/SUM[12] ) );
  XNOR2_X1 U5643 ( .A(n4207), .B(n4070), .ZN(n5003) );
  AOI22_X1 U5644 ( .A1(n3898), .A2(\dp/id_exe_regs/b_mult_reg/q[27] ), .B1(
        n3956), .B2(\dp/id_exe_regs/b_mult_reg/q[29] ), .ZN(n6961) );
  NAND2_X1 U5645 ( .A1(n5213), .A2(\dp/ids/rp2[28] ), .ZN(n6962) );
  AOI22_X1 U5646 ( .A1(n3898), .A2(\dp/id_exe_regs/b_mult_reg/q[26] ), .B1(
        n3947), .B2(\dp/id_exe_regs/b_mult_reg/q[28] ), .ZN(n6924) );
  NAND2_X1 U5647 ( .A1(n5214), .A2(\dp/ids/rp2[27] ), .ZN(n6925) );
  NAND2_X1 U5648 ( .A1(n6923), .A2(n6928), .ZN(n6963) );
  OAI21_X1 U5649 ( .B1(n7147), .B2(b_selector_id), .A(n6922), .ZN(n6928) );
  INV_X1 U5650 ( .A(n6980), .ZN(n6922) );
  NAND2_X1 U5651 ( .A1(n6921), .A2(is_signed_id), .ZN(n7147) );
  NOR2_X1 U5652 ( .A1(n4360), .A2(sign_ext_sel_id), .ZN(n6921) );
  OAI22_X1 U5653 ( .A1(n6621), .A2(n5196), .B1(n6620), .B2(n4808), .ZN(n2831)
         );
  XNOR2_X1 U5654 ( .A(n4918), .B(n6619), .ZN(n6621) );
  NOR2_X1 U5655 ( .A1(n6618), .A2(n6617), .ZN(n6619) );
  INV_X1 U5656 ( .A(n6616), .ZN(n6618) );
  AOI21_X1 U5657 ( .B1(n6714), .B2(n4920), .A(n4919), .ZN(n4918) );
  OAI21_X1 U5658 ( .B1(n6646), .B2(n6607), .A(n6606), .ZN(n6614) );
  INV_X1 U5659 ( .A(n6605), .ZN(n6606) );
  AND2_X1 U5660 ( .A1(n6612), .A2(n6615), .ZN(n4920) );
  NOR2_X1 U5661 ( .A1(n6642), .A2(n6607), .ZN(n6612) );
  OAI22_X1 U5662 ( .A1(n6698), .A2(n7062), .B1(n7434), .B2(n3938), .ZN(n2790)
         );
  XNOR2_X1 U5663 ( .A(n6697), .B(n6696), .ZN(n6698) );
  NOR2_X1 U5664 ( .A1(n6703), .A2(n6700), .ZN(n6696) );
  INV_X1 U5665 ( .A(n6699), .ZN(n6695) );
  OAI22_X1 U5666 ( .A1(n5198), .A2(n6577), .B1(n4406), .B2(n4808), .ZN(n2837)
         );
  INV_X1 U5667 ( .A(n7098), .ZN(n4808) );
  XNOR2_X1 U5668 ( .A(n6576), .B(n6575), .ZN(n6577) );
  NOR2_X1 U5669 ( .A1(n6574), .A2(n6573), .ZN(n6575) );
  INV_X1 U5670 ( .A(n6572), .ZN(n6574) );
  NAND2_X1 U5671 ( .A1(n6560), .A2(n6562), .ZN(n6578) );
  INV_X1 U5672 ( .A(n6534), .ZN(n6560) );
  INV_X1 U5673 ( .A(n6571), .ZN(n6567) );
  INV_X1 U5674 ( .A(n6581), .ZN(n6570) );
  AOI21_X1 U5675 ( .B1(n6563), .B2(n6562), .A(n6561), .ZN(n6581) );
  OAI22_X1 U5676 ( .A1(n7063), .A2(n5198), .B1(n4583), .B2(n5199), .ZN(n2819)
         );
  OAI22_X1 U5677 ( .A1(n6509), .A2(n5196), .B1(n4473), .B2(n5199), .ZN(n2845)
         );
  OAI22_X1 U5678 ( .A1(n5563), .A2(n5561), .B1(n3935), .B2(n4542), .ZN(
        \ctrl_u/n547 ) );
  NAND2_X1 U5679 ( .A1(n5627), .A2(n5560), .ZN(n5561) );
  AND2_X1 U5680 ( .A1(n3929), .A2(n5038), .ZN(n4844) );
  OAI22_X1 U5681 ( .A1(n5557), .A2(n5556), .B1(n3935), .B2(n4540), .ZN(
        \ctrl_u/n545 ) );
  INV_X1 U5682 ( .A(n5562), .ZN(n5556) );
  AOI22_X1 U5683 ( .A1(n3894), .A2(\dp/ifs/pc_btb[29] ), .B1(n5193), .B2(
        btb_cache_read_address[29]), .ZN(n6184) );
  OAI21_X1 U5684 ( .B1(n6162), .B2(n7069), .A(n6158), .ZN(n6160) );
  NAND2_X1 U5685 ( .A1(n6162), .A2(n3952), .ZN(n6158) );
  OAI22_X1 U5686 ( .A1(n6660), .A2(n5196), .B1(n4385), .B2(n5199), .ZN(n2827)
         );
  OAI22_X1 U5687 ( .A1(n6641), .A2(n5196), .B1(n4382), .B2(n5199), .ZN(n2829)
         );
  OAI211_X1 U5688 ( .C1(n3935), .C2(n4580), .A(n5570), .B(n5547), .ZN(
        \ctrl_u/n522 ) );
  OAI21_X1 U5689 ( .B1(n5496), .B2(n5502), .A(n5495), .ZN(n4856) );
  NOR2_X1 U5690 ( .A1(n5604), .A2(n5587), .ZN(n5495) );
  OAI211_X1 U5691 ( .C1(n3873), .C2(\intadd_2/B[14] ), .A(n6388), .B(n6387), 
        .ZN(n2542) );
  AOI22_X1 U5692 ( .A1(n3931), .A2(\dp/ifs/pc_btb[15] ), .B1(n7108), .B2(
        btb_cache_read_address[15]), .ZN(n6387) );
  NOR2_X1 U5693 ( .A1(n6386), .A2(n4908), .ZN(n6388) );
  NAND2_X1 U5694 ( .A1(n4911), .A2(n4909), .ZN(n4908) );
  NAND2_X1 U5695 ( .A1(n3883), .A2(n4910), .ZN(n4909) );
  AOI21_X1 U5696 ( .B1(n5766), .B2(n7076), .A(n5765), .ZN(n7438) );
  OAI211_X1 U5697 ( .C1(\intadd_1/SUM[16] ), .C2(n7066), .A(n5764), .B(n5763), 
        .ZN(n5765) );
  NAND2_X1 U5698 ( .A1(n5111), .A2(n3952), .ZN(n5761) );
  INV_X1 U5699 ( .A(n5760), .ZN(n5111) );
  NAND2_X1 U5700 ( .A1(\dp/exs/alu_unit/shifter_out[17] ), .A2(n3954), .ZN(
        n5764) );
  XNOR2_X1 U5701 ( .A(n5956), .B(n5955), .ZN(n5759) );
  AOI21_X1 U5702 ( .B1(n5758), .B2(n5103), .A(n4106), .ZN(n5100) );
  NAND2_X1 U5703 ( .A1(n4784), .A2(n4787), .ZN(n5758) );
  NAND2_X1 U5704 ( .A1(n5945), .A2(n4814), .ZN(n4784) );
  NAND2_X1 U5705 ( .A1(n4993), .A2(n4992), .ZN(n5931) );
  NAND2_X1 U5706 ( .A1(n3936), .A2(\dp/pc_plus4_out_if_int[15] ), .ZN(n4911)
         );
  NOR2_X1 U5707 ( .A1(n3879), .A2(\intadd_2/SUM[14] ), .ZN(n6386) );
  OAI21_X1 U5708 ( .B1(n6482), .B2(n5198), .A(n4810), .ZN(n2849) );
  NAND2_X1 U5709 ( .A1(n7098), .A2(\dp/a_neg_mult_id_exe_int[33] ), .ZN(n4810)
         );
  INV_X1 U5710 ( .A(n7181), .ZN(n280) );
  AOI22_X1 U5711 ( .A1(n5133), .A2(rs_id[1]), .B1(n5180), .B2(instr_if[22]), 
        .ZN(n7181) );
  NAND2_X1 U5712 ( .A1(n3928), .A2(\dp/pc_plus4_out_if_int[27] ), .ZN(n6403)
         );
  AOI22_X1 U5713 ( .A1(n3895), .A2(\dp/ifs/pc_btb[27] ), .B1(n5193), .B2(
        btb_cache_read_address[27]), .ZN(n6404) );
  OAI22_X1 U5714 ( .A1(n6509), .A2(n7062), .B1(n4172), .B2(n7439), .ZN(n2813)
         );
  XNOR2_X1 U5715 ( .A(n6508), .B(n6507), .ZN(n6509) );
  NOR2_X1 U5716 ( .A1(n6506), .A2(n6505), .ZN(n6507) );
  INV_X1 U5717 ( .A(n6501), .ZN(n6504) );
  OAI22_X1 U5718 ( .A1(n7063), .A2(n7062), .B1(n681), .B2(n3942), .ZN(n2787)
         );
  XNOR2_X1 U5719 ( .A(n6332), .B(n6331), .ZN(n7063) );
  OAI211_X1 U5720 ( .C1(n681), .C2(n3930), .A(n6325), .B(n6324), .ZN(n6330) );
  NAND2_X1 U5721 ( .A1(n3943), .A2(\dp/a_neg_mult_id_exe_int[62] ), .ZN(n6324)
         );
  OR2_X1 U5722 ( .A1(n6699), .A2(n6319), .ZN(n6711) );
  NAND2_X1 U5723 ( .A1(n6693), .A2(n6690), .ZN(n6699) );
  NOR2_X1 U5724 ( .A1(n6684), .A2(n6318), .ZN(n6693) );
  NAND2_X1 U5725 ( .A1(n6622), .A2(n6317), .ZN(n6684) );
  NOR2_X1 U5726 ( .A1(n6305), .A2(n6304), .ZN(n6715) );
  NOR2_X1 U5727 ( .A1(n6302), .A2(n6301), .ZN(n6706) );
  NOR2_X1 U5728 ( .A1(n6300), .A2(n6299), .ZN(n6703) );
  NAND2_X1 U5729 ( .A1(n6303), .A2(n6705), .ZN(n6319) );
  INV_X1 U5730 ( .A(n6700), .ZN(n6705) );
  AND2_X1 U5731 ( .A1(n6300), .A2(n6299), .ZN(n6700) );
  INV_X1 U5732 ( .A(n6707), .ZN(n6303) );
  AND2_X1 U5733 ( .A1(n6302), .A2(n6301), .ZN(n6707) );
  NAND2_X1 U5734 ( .A1(n6297), .A2(n6691), .ZN(n6704) );
  NAND2_X1 U5735 ( .A1(n6692), .A2(n6690), .ZN(n6297) );
  NAND2_X1 U5736 ( .A1(n6295), .A2(n6296), .ZN(n6690) );
  NAND2_X1 U5737 ( .A1(n6294), .A2(n6685), .ZN(n6692) );
  NAND2_X1 U5738 ( .A1(n6682), .A2(n6686), .ZN(n6294) );
  INV_X1 U5739 ( .A(n6318), .ZN(n6686) );
  AND2_X1 U5740 ( .A1(n6292), .A2(n6293), .ZN(n6318) );
  NOR2_X1 U5741 ( .A1(n6645), .A2(n6282), .ZN(n6317) );
  NAND2_X1 U5742 ( .A1(n6287), .A2(n6664), .ZN(n6282) );
  AND2_X1 U5743 ( .A1(n6676), .A2(n6675), .ZN(n6287) );
  INV_X1 U5744 ( .A(n6716), .ZN(n6321) );
  AND2_X1 U5745 ( .A1(n6305), .A2(n6304), .ZN(n6716) );
  NOR3_X1 U5746 ( .A1(n5576), .A2(n5509), .A3(n5508), .ZN(n5568) );
  OAI21_X1 U5747 ( .B1(n5507), .B2(n5506), .A(n5505), .ZN(n5508) );
  NAND2_X1 U5748 ( .A1(n5553), .A2(n5558), .ZN(n5505) );
  NOR2_X1 U5749 ( .A1(instr_if[28]), .A2(n5490), .ZN(n5558) );
  AOI21_X1 U5750 ( .B1(instr_if[30]), .B2(n5560), .A(n5588), .ZN(n5507) );
  OAI211_X1 U5751 ( .C1(n5514), .C2(n5587), .A(n5511), .B(n5625), .ZN(n5509)
         );
  NAND2_X1 U5752 ( .A1(n5552), .A2(n5644), .ZN(n5511) );
  OAI211_X1 U5753 ( .C1(n4361), .C2(n7165), .A(n7142), .B(n7168), .ZN(n3067)
         );
  AOI22_X1 U5754 ( .A1(n7164), .A2(rt_id[0]), .B1(n7166), .B2(rd_idexe[0]), 
        .ZN(n7142) );
  OAI211_X1 U5755 ( .C1(n4363), .C2(n7165), .A(n7144), .B(n7168), .ZN(n3065)
         );
  AOI22_X1 U5756 ( .A1(n7164), .A2(rt_id[2]), .B1(n7166), .B2(rd_idexe[2]), 
        .ZN(n7144) );
  OAI211_X1 U5757 ( .C1(n4364), .C2(n7165), .A(n7145), .B(n7168), .ZN(n3064)
         );
  AOI22_X1 U5758 ( .A1(n7164), .A2(rt_id[3]), .B1(n7166), .B2(rd_idexe[3]), 
        .ZN(n7145) );
  OAI211_X1 U5759 ( .C1(n4362), .C2(n7165), .A(n7143), .B(n7168), .ZN(n3066)
         );
  AOI22_X1 U5760 ( .A1(n7164), .A2(rt_id[1]), .B1(n7166), .B2(rd_idexe[1]), 
        .ZN(n7143) );
  OAI22_X1 U5761 ( .A1(n6660), .A2(n7062), .B1(n4186), .B2(n3942), .ZN(n2795)
         );
  XNOR2_X1 U5762 ( .A(n6659), .B(n6658), .ZN(n6660) );
  NOR2_X1 U5763 ( .A1(n6657), .A2(n6656), .ZN(n6658) );
  INV_X1 U5764 ( .A(n6655), .ZN(n6657) );
  INV_X1 U5765 ( .A(n6661), .ZN(n6650) );
  OAI22_X1 U5766 ( .A1(n6681), .A2(n7062), .B1(n4177), .B2(n3938), .ZN(n2793)
         );
  XNOR2_X1 U5767 ( .A(n6680), .B(n6679), .ZN(n6681) );
  NOR2_X1 U5768 ( .A1(n6678), .A2(n6677), .ZN(n6679) );
  NOR2_X1 U5769 ( .A1(n6291), .A2(n6290), .ZN(n6677) );
  INV_X1 U5770 ( .A(n6676), .ZN(n6678) );
  NAND2_X1 U5771 ( .A1(n6291), .A2(n6290), .ZN(n6676) );
  NAND2_X1 U5772 ( .A1(n6661), .A2(n6664), .ZN(n6670) );
  INV_X1 U5773 ( .A(n6675), .ZN(n6671) );
  NOR2_X1 U5774 ( .A1(n6289), .A2(n6288), .ZN(n6673) );
  INV_X1 U5775 ( .A(n6669), .ZN(n6674) );
  AOI21_X1 U5776 ( .B1(n6665), .B2(n6664), .A(n6663), .ZN(n6669) );
  INV_X1 U5777 ( .A(n6662), .ZN(n6663) );
  AOI21_X1 U5778 ( .B1(n6653), .B2(n6655), .A(n6656), .ZN(n6662) );
  NOR2_X1 U5779 ( .A1(n6286), .A2(n6285), .ZN(n6656) );
  AND2_X1 U5780 ( .A1(n6654), .A2(n6655), .ZN(n6664) );
  NAND2_X1 U5781 ( .A1(n6286), .A2(n6285), .ZN(n6655) );
  NAND2_X1 U5782 ( .A1(n6289), .A2(n6288), .ZN(n6675) );
  OAI21_X1 U5783 ( .B1(n6596), .B2(n5197), .A(n4811), .ZN(n2834) );
  NAND2_X1 U5784 ( .A1(n7098), .A2(\dp/a_neg_mult_id_exe_int[48] ), .ZN(n4811)
         );
  OAI22_X1 U5785 ( .A1(n6641), .A2(n7062), .B1(n4176), .B2(n3942), .ZN(n2797)
         );
  XNOR2_X1 U5786 ( .A(n6640), .B(n6639), .ZN(n6641) );
  NOR2_X1 U5787 ( .A1(n6638), .A2(n6637), .ZN(n6639) );
  INV_X1 U5788 ( .A(n6636), .ZN(n6638) );
  NAND2_X1 U5789 ( .A1(n6622), .A2(n6624), .ZN(n6630) );
  INV_X1 U5790 ( .A(n6635), .ZN(n6631) );
  INV_X1 U5791 ( .A(n6629), .ZN(n6634) );
  AOI21_X1 U5792 ( .B1(n6625), .B2(n6624), .A(n6623), .ZN(n6629) );
  OAI21_X1 U5793 ( .B1(n6649), .B2(n5196), .A(n4812), .ZN(n2828) );
  NAND2_X1 U5794 ( .A1(n7098), .A2(\dp/a_neg_mult_id_exe_int[54] ), .ZN(n4812)
         );
  NAND2_X1 U5795 ( .A1(n4806), .A2(n4805), .ZN(\ctrl_u/n512 ) );
  NAND2_X1 U5796 ( .A1(n5181), .A2(n4481), .ZN(n4805) );
  INV_X1 U5797 ( .A(n4807), .ZN(n4806) );
  OAI22_X1 U5798 ( .A1(n5584), .A2(n5583), .B1(n3927), .B2(n5582), .ZN(n4807)
         );
  AOI211_X1 U5799 ( .C1(instr_if[3]), .C2(n5580), .A(n5579), .B(n5578), .ZN(
        n5582) );
  OAI211_X1 U5800 ( .C1(n5596), .C2(n5519), .A(n5624), .B(n5531), .ZN(n5578)
         );
  NOR2_X1 U5801 ( .A1(n5595), .A2(n5596), .ZN(n5498) );
  INV_X1 U5802 ( .A(n5577), .ZN(n5580) );
  NOR3_X1 U5803 ( .A1(n5576), .A2(n5575), .A3(n5574), .ZN(n5583) );
  OAI211_X1 U5804 ( .C1(instr_if[30]), .C2(n5633), .A(n5573), .B(n5572), .ZN(
        n5574) );
  NAND2_X1 U5805 ( .A1(n5553), .A2(n5646), .ZN(n5572) );
  NOR2_X1 U5806 ( .A1(instr_if[27]), .A2(instr_if[29]), .ZN(n5646) );
  NAND2_X1 U5807 ( .A1(n5649), .A2(n7276), .ZN(n5573) );
  OAI211_X1 U5808 ( .C1(n7276), .C2(n5651), .A(n5512), .B(n5625), .ZN(n5575)
         );
  NAND2_X1 U5809 ( .A1(n5504), .A2(n5650), .ZN(n5625) );
  INV_X1 U5810 ( .A(n5491), .ZN(n5650) );
  AOI21_X1 U5811 ( .B1(n5506), .B2(n5503), .A(n7275), .ZN(n5576) );
  NAND2_X1 U5812 ( .A1(n5496), .A2(n5638), .ZN(n5513) );
  NOR3_X1 U5813 ( .A1(n3886), .A2(n6599), .A3(n6642), .ZN(n6600) );
  NOR3_X1 U5814 ( .A1(n3872), .A2(n6535), .A3(n6534), .ZN(n6536) );
  INV_X1 U5815 ( .A(n6538), .ZN(n6535) );
  NAND2_X1 U5816 ( .A1(n6887), .A2(n6886), .ZN(n2945) );
  NAND2_X1 U5817 ( .A1(n5202), .A2(n6885), .ZN(n6886) );
  INV_X1 U5818 ( .A(n6889), .ZN(n6885) );
  NAND2_X1 U5819 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[1] ), .ZN(n6887) );
  NAND2_X1 U5820 ( .A1(n6871), .A2(n6870), .ZN(n2941) );
  NAND2_X1 U5821 ( .A1(n5202), .A2(n6869), .ZN(n6870) );
  INV_X1 U5822 ( .A(n6873), .ZN(n6869) );
  NAND2_X1 U5823 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[5] ), .ZN(n6871) );
  NAND2_X1 U5824 ( .A1(n6877), .A2(n6876), .ZN(n2942) );
  NAND2_X1 U5825 ( .A1(n5200), .A2(n6875), .ZN(n6876) );
  INV_X1 U5826 ( .A(n6879), .ZN(n6875) );
  NAND2_X1 U5827 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[4] ), .ZN(n6877) );
  NAND2_X1 U5828 ( .A1(n6892), .A2(n6891), .ZN(n2946) );
  NAND2_X1 U5829 ( .A1(n7056), .A2(n6890), .ZN(n6891) );
  INV_X1 U5830 ( .A(n6894), .ZN(n6890) );
  NAND2_X1 U5831 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[0] ), .ZN(n6892) );
  NAND2_X1 U5832 ( .A1(n6809), .A2(n6808), .ZN(n2924) );
  NAND2_X1 U5833 ( .A1(n5202), .A2(n6807), .ZN(n6808) );
  INV_X1 U5834 ( .A(n6811), .ZN(n6807) );
  NAND2_X1 U5835 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[22] ), .ZN(n6809) );
  NAND2_X1 U5836 ( .A1(n6798), .A2(n6797), .ZN(n2922) );
  NAND2_X1 U5837 ( .A1(n5202), .A2(n6796), .ZN(n6797) );
  INV_X1 U5838 ( .A(n6800), .ZN(n6796) );
  NAND2_X1 U5839 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[24] ), .ZN(n6798) );
  NAND2_X1 U5840 ( .A1(n6780), .A2(n6779), .ZN(n2919) );
  NAND2_X1 U5841 ( .A1(n5201), .A2(n6778), .ZN(n6779) );
  INV_X1 U5842 ( .A(n6782), .ZN(n6778) );
  NAND2_X1 U5843 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[27] ), .ZN(n6780) );
  NAND2_X1 U5844 ( .A1(n6804), .A2(n6803), .ZN(n2923) );
  NAND2_X1 U5845 ( .A1(n5200), .A2(n6802), .ZN(n6803) );
  INV_X1 U5846 ( .A(n6806), .ZN(n6802) );
  NAND2_X1 U5847 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[23] ), .ZN(n6804) );
  NAND2_X1 U5848 ( .A1(n6814), .A2(n6813), .ZN(n2925) );
  NAND2_X1 U5849 ( .A1(n5201), .A2(n6812), .ZN(n6813) );
  INV_X1 U5850 ( .A(n6816), .ZN(n6812) );
  NAND2_X1 U5851 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[21] ), .ZN(n6814) );
  NAND2_X1 U5852 ( .A1(n6830), .A2(n6829), .ZN(n2928) );
  NAND2_X1 U5853 ( .A1(n5201), .A2(n6828), .ZN(n6829) );
  INV_X1 U5854 ( .A(n6832), .ZN(n6828) );
  NAND2_X1 U5855 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[18] ), .ZN(n6830) );
  NAND2_X1 U5856 ( .A1(n6774), .A2(n6773), .ZN(n2918) );
  NAND2_X1 U5857 ( .A1(n5201), .A2(n6772), .ZN(n6773) );
  INV_X1 U5858 ( .A(n6776), .ZN(n6772) );
  NAND2_X1 U5859 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[28] ), .ZN(n6774) );
  NAND2_X1 U5860 ( .A1(n6762), .A2(n6761), .ZN(n2916) );
  NAND2_X1 U5861 ( .A1(n5202), .A2(n6760), .ZN(n6761) );
  INV_X1 U5862 ( .A(n6764), .ZN(n6760) );
  NAND2_X1 U5863 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[30] ), .ZN(n6762) );
  NAND2_X1 U5864 ( .A1(n6768), .A2(n6767), .ZN(n2917) );
  NAND2_X1 U5865 ( .A1(n5200), .A2(n6766), .ZN(n6767) );
  INV_X1 U5866 ( .A(n6770), .ZN(n6766) );
  NAND2_X1 U5867 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[29] ), .ZN(n6768) );
  NAND2_X1 U5868 ( .A1(n6824), .A2(n6823), .ZN(n2927) );
  NAND2_X1 U5869 ( .A1(n7056), .A2(n6822), .ZN(n6823) );
  INV_X1 U5870 ( .A(n6826), .ZN(n6822) );
  NAND2_X1 U5871 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[19] ), .ZN(n6824) );
  NAND2_X1 U5872 ( .A1(n6792), .A2(n6791), .ZN(n2921) );
  NAND2_X1 U5873 ( .A1(n7056), .A2(n6790), .ZN(n6791) );
  INV_X1 U5874 ( .A(n6794), .ZN(n6790) );
  NAND2_X1 U5875 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[25] ), .ZN(n6792) );
  NOR2_X1 U5876 ( .A1(n6599), .A2(n6601), .ZN(n6594) );
  INV_X1 U5877 ( .A(n6602), .ZN(n6599) );
  NOR2_X1 U5878 ( .A1(n6651), .A2(n6653), .ZN(n6647) );
  NOR2_X1 U5879 ( .A1(n6284), .A2(n6283), .ZN(n6653) );
  INV_X1 U5880 ( .A(n6654), .ZN(n6651) );
  NAND2_X1 U5881 ( .A1(n6284), .A2(n6283), .ZN(n6654) );
  OAI21_X1 U5882 ( .B1(n6646), .B2(n6645), .A(n6644), .ZN(n6665) );
  INV_X1 U5883 ( .A(n6643), .ZN(n6644) );
  NAND2_X1 U5884 ( .A1(n6281), .A2(n6280), .ZN(n6643) );
  AOI21_X1 U5885 ( .B1(n6633), .B2(n6636), .A(n6637), .ZN(n6280) );
  NOR2_X1 U5886 ( .A1(n6279), .A2(n6278), .ZN(n6637) );
  NOR2_X1 U5887 ( .A1(n6277), .A2(n6276), .ZN(n6633) );
  NAND2_X1 U5888 ( .A1(n6623), .A2(n6275), .ZN(n6281) );
  NOR2_X1 U5889 ( .A1(n6274), .A2(n6273), .ZN(n6617) );
  NOR2_X1 U5890 ( .A1(n6272), .A2(n6271), .ZN(n6613) );
  NAND2_X1 U5891 ( .A1(n6269), .A2(n6598), .ZN(n6605) );
  NAND2_X1 U5892 ( .A1(n6601), .A2(n6597), .ZN(n6269) );
  NOR2_X1 U5893 ( .A1(n6266), .A2(n6265), .ZN(n6601) );
  INV_X1 U5894 ( .A(n6625), .ZN(n6646) );
  NAND2_X1 U5895 ( .A1(n6259), .A2(n6258), .ZN(n6625) );
  AOI21_X1 U5896 ( .B1(n6257), .B2(n6561), .A(n6256), .ZN(n6258) );
  OAI21_X1 U5897 ( .B1(n6579), .B2(n6255), .A(n6254), .ZN(n6256) );
  AOI21_X1 U5898 ( .B1(n6587), .B2(n6590), .A(n6591), .ZN(n6254) );
  NOR2_X1 U5899 ( .A1(n6253), .A2(n6252), .ZN(n6591) );
  NOR2_X1 U5900 ( .A1(n6251), .A2(n6250), .ZN(n6587) );
  AOI21_X1 U5901 ( .B1(n6569), .B2(n6572), .A(n6573), .ZN(n6579) );
  NOR2_X1 U5902 ( .A1(n6249), .A2(n6248), .ZN(n6573) );
  NOR2_X1 U5903 ( .A1(n6247), .A2(n6246), .ZN(n6569) );
  NOR2_X1 U5904 ( .A1(n6245), .A2(n6244), .ZN(n6555) );
  NOR2_X1 U5905 ( .A1(n6243), .A2(n6242), .ZN(n6551) );
  NAND2_X1 U5906 ( .A1(n6240), .A2(n6533), .ZN(n6542) );
  NAND2_X1 U5907 ( .A1(n6537), .A2(n6532), .ZN(n6240) );
  NOR2_X1 U5908 ( .A1(n6237), .A2(n6236), .ZN(n6537) );
  NAND2_X1 U5909 ( .A1(n6563), .A2(n6235), .ZN(n6259) );
  INV_X1 U5910 ( .A(n6316), .ZN(n6235) );
  NOR2_X1 U5911 ( .A1(n6642), .A2(n6645), .ZN(n6661) );
  NAND2_X1 U5912 ( .A1(n6624), .A2(n6275), .ZN(n6645) );
  AND2_X1 U5913 ( .A1(n6635), .A2(n6636), .ZN(n6275) );
  NAND2_X1 U5914 ( .A1(n6279), .A2(n6278), .ZN(n6636) );
  NAND2_X1 U5915 ( .A1(n6277), .A2(n6276), .ZN(n6635) );
  NOR2_X1 U5916 ( .A1(n6607), .A2(n6270), .ZN(n6624) );
  NAND2_X1 U5917 ( .A1(n6615), .A2(n6616), .ZN(n6270) );
  NAND2_X1 U5918 ( .A1(n6274), .A2(n6273), .ZN(n6616) );
  NAND2_X1 U5919 ( .A1(n6272), .A2(n6271), .ZN(n6615) );
  NAND4_X1 U5920 ( .A1(n6264), .A2(n6263), .A3(n6262), .A4(n6261), .ZN(n6272)
         );
  NAND2_X1 U5921 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[50] ), .A2(n3946), 
        .ZN(n6261) );
  NAND2_X1 U5922 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[49] ), .A2(n5189), .ZN(
        n6262) );
  NAND2_X1 U5923 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[49] ), .A2(n6326), 
        .ZN(n6263) );
  AOI21_X1 U5924 ( .B1(\dp/exs/alu_unit/mult/a_shiftn[50] ), .B2(n3945), .A(
        n6260), .ZN(n6264) );
  NOR2_X1 U5925 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[50] ), .ZN(n6260) );
  NAND2_X1 U5926 ( .A1(n6602), .A2(n6597), .ZN(n6607) );
  NAND2_X1 U5927 ( .A1(n6267), .A2(n6268), .ZN(n6597) );
  NAND2_X1 U5928 ( .A1(n6266), .A2(n6265), .ZN(n6602) );
  INV_X1 U5929 ( .A(n6622), .ZN(n6642) );
  NOR2_X1 U5930 ( .A1(n6534), .A2(n6316), .ZN(n6622) );
  NAND2_X1 U5931 ( .A1(n6562), .A2(n6257), .ZN(n6316) );
  NOR2_X1 U5932 ( .A1(n6580), .A2(n6255), .ZN(n6257) );
  NAND2_X1 U5933 ( .A1(n6589), .A2(n6590), .ZN(n6255) );
  NAND2_X1 U5934 ( .A1(n6253), .A2(n6252), .ZN(n6590) );
  NAND2_X1 U5935 ( .A1(n6251), .A2(n6250), .ZN(n6589) );
  NAND2_X1 U5936 ( .A1(n6571), .A2(n6572), .ZN(n6580) );
  NAND2_X1 U5937 ( .A1(n6249), .A2(n6248), .ZN(n6572) );
  NAND4_X1 U5938 ( .A1(n6234), .A2(n6233), .A3(n6232), .A4(n6231), .ZN(n6249)
         );
  NAND2_X1 U5939 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[44] ), .A2(n5189), .ZN(
        n6231) );
  NAND2_X1 U5940 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[44] ), .A2(n5154), 
        .ZN(n6232) );
  NAND2_X1 U5941 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[45] ), .A2(n3946), 
        .ZN(n6233) );
  AOI21_X1 U5942 ( .B1(\dp/exs/alu_unit/mult/a_shiftn[45] ), .B2(n3945), .A(
        n6230), .ZN(n6234) );
  NOR2_X1 U5943 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[45] ), .ZN(n6230) );
  NAND2_X1 U5944 ( .A1(n6247), .A2(n6246), .ZN(n6571) );
  NAND4_X1 U5945 ( .A1(n6229), .A2(n6228), .A3(n6227), .A4(n6226), .ZN(n6247)
         );
  NAND2_X1 U5946 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[44] ), .A2(n3946), 
        .ZN(n6226) );
  NAND2_X1 U5947 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[43] ), .A2(n5189), .ZN(
        n6227) );
  NAND2_X1 U5948 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[43] ), .A2(n5154), 
        .ZN(n6228) );
  AOI21_X1 U5949 ( .B1(\dp/exs/alu_unit/mult/a_shiftn[44] ), .B2(n3945), .A(
        n6225), .ZN(n6229) );
  NOR2_X1 U5950 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[44] ), .ZN(n6225) );
  NOR2_X1 U5951 ( .A1(n6241), .A2(n6541), .ZN(n6562) );
  NAND2_X1 U5952 ( .A1(n6538), .A2(n6532), .ZN(n6541) );
  NAND2_X1 U5953 ( .A1(n6238), .A2(n6239), .ZN(n6532) );
  NAND4_X1 U5954 ( .A1(n6224), .A2(n6223), .A3(n6222), .A4(n6221), .ZN(n6238)
         );
  NAND2_X1 U5955 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[40] ), .A2(n5154), 
        .ZN(n6221) );
  NAND2_X1 U5956 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[40] ), .A2(n6298), .ZN(
        n6222) );
  NAND2_X1 U5957 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[41] ), .A2(n3945), .ZN(
        n6223) );
  AOI21_X1 U5958 ( .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[41] ), .B2(n5188), 
        .A(n6220), .ZN(n6224) );
  NOR2_X1 U5959 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[41] ), .ZN(n6220) );
  NAND2_X1 U5960 ( .A1(n6237), .A2(n6236), .ZN(n6538) );
  NAND2_X1 U5961 ( .A1(n6554), .A2(n6553), .ZN(n6241) );
  NAND2_X1 U5962 ( .A1(n6243), .A2(n6242), .ZN(n6553) );
  NAND2_X1 U5963 ( .A1(n6245), .A2(n6244), .ZN(n6554) );
  NAND2_X1 U5964 ( .A1(n6513), .A2(n6219), .ZN(n6315) );
  AND2_X1 U5965 ( .A1(n6518), .A2(n6526), .ZN(n6219) );
  AOI22_X1 U5966 ( .A1(n5134), .A2(\dp/imm_id_int[4] ), .B1(n5179), .B2(
        instr_if[4]), .ZN(n1638) );
  AOI22_X1 U5967 ( .A1(n5134), .A2(\dp/imm_id_int[5] ), .B1(n5179), .B2(
        instr_if[5]), .ZN(n1637) );
  AOI22_X1 U5968 ( .A1(n5133), .A2(\dp/imm_id_int[12] ), .B1(n5179), .B2(
        instr_if[12]), .ZN(n1630) );
  INV_X1 U5969 ( .A(n3924), .ZN(n5654) );
  OAI21_X1 U5970 ( .B1(n6528), .B2(n5196), .A(n4813), .ZN(n2843) );
  NAND2_X1 U5971 ( .A1(n7098), .A2(\dp/a_neg_mult_id_exe_int[39] ), .ZN(n4813)
         );
  NOR3_X1 U5972 ( .A1(n3886), .A2(n6522), .A3(n6521), .ZN(n6523) );
  NAND2_X1 U5973 ( .A1(n6511), .A2(n6513), .ZN(n6521) );
  INV_X1 U5974 ( .A(n6510), .ZN(n6511) );
  NAND2_X1 U5975 ( .A1(n6486), .A2(n6314), .ZN(n6510) );
  NAND2_X1 U5976 ( .A1(n6313), .A2(n6312), .ZN(n6480) );
  INV_X1 U5977 ( .A(n6526), .ZN(n6522) );
  AOI21_X1 U5978 ( .B1(n6146), .B2(n6306), .A(n6307), .ZN(n4869) );
  NAND2_X1 U5979 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[30] ), .A2(n5189), .ZN(
        n6152) );
  NAND2_X1 U5980 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[31] ), .A2(n3946), 
        .ZN(n6153) );
  NAND2_X1 U5981 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[31] ), .A2(n3945), .ZN(
        n6154) );
  AOI21_X1 U5982 ( .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[30] ), .B2(n5154), 
        .A(n6151), .ZN(n6155) );
  NOR2_X1 U5983 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[31] ), .ZN(n6151) );
  OAI21_X1 U5984 ( .B1(n6145), .B2(n6144), .A(n6143), .ZN(n6146) );
  AOI22_X1 U5985 ( .A1(n6142), .A2(n6141), .B1(n6140), .B2(n6139), .ZN(n6143)
         );
  NAND2_X1 U5986 ( .A1(n6150), .A2(n6149), .ZN(n6306) );
  AOI22_X1 U5987 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[31] ), .B1(n5156), 
        .B2(\dp/mul_feedback_exe_mem_int[31] ), .ZN(n6149) );
  AOI22_X1 U5988 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[30] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[31] ), .ZN(n6150) );
  OAI21_X1 U5989 ( .B1(n6138), .B2(n6144), .A(n6145), .ZN(n6147) );
  NAND2_X1 U5990 ( .A1(n6137), .A2(n6136), .ZN(n6145) );
  INV_X1 U5991 ( .A(n6135), .ZN(n6144) );
  INV_X1 U5992 ( .A(n6137), .ZN(n6138) );
  NOR2_X1 U5993 ( .A1(n6134), .A2(n6133), .ZN(n6142) );
  NOR2_X1 U5994 ( .A1(n6139), .A2(n6140), .ZN(n6134) );
  NOR2_X1 U5995 ( .A1(n6216), .A2(n6215), .ZN(n6524) );
  INV_X1 U5996 ( .A(n6520), .ZN(n6525) );
  AOI21_X1 U5997 ( .B1(n6514), .B2(n6513), .A(n6512), .ZN(n6520) );
  OAI21_X1 U5998 ( .B1(n6497), .B2(n6506), .A(n6214), .ZN(n6512) );
  INV_X1 U5999 ( .A(n6505), .ZN(n6214) );
  NOR2_X1 U6000 ( .A1(n6213), .A2(n6212), .ZN(n6505) );
  INV_X1 U6001 ( .A(n6503), .ZN(n6497) );
  NOR2_X1 U6002 ( .A1(n6211), .A2(n6210), .ZN(n6503) );
  NOR2_X1 U6003 ( .A1(n6501), .A2(n6506), .ZN(n6513) );
  AND2_X1 U6004 ( .A1(n6213), .A2(n6212), .ZN(n6506) );
  AND2_X1 U6005 ( .A1(n6211), .A2(n6210), .ZN(n6501) );
  NAND2_X1 U6006 ( .A1(n6204), .A2(n6203), .ZN(n6514) );
  AOI21_X1 U6007 ( .B1(n6489), .B2(n6492), .A(n6493), .ZN(n6203) );
  NOR2_X1 U6008 ( .A1(n6202), .A2(n6201), .ZN(n6493) );
  NOR2_X1 U6009 ( .A1(n6200), .A2(n6199), .ZN(n6489) );
  NAND2_X1 U6010 ( .A1(n6490), .A2(n6314), .ZN(n6204) );
  AND2_X1 U6011 ( .A1(n6491), .A2(n6492), .ZN(n6314) );
  NAND2_X1 U6012 ( .A1(n6202), .A2(n6201), .ZN(n6492) );
  NAND2_X1 U6013 ( .A1(n6200), .A2(n6199), .ZN(n6491) );
  NAND2_X1 U6014 ( .A1(n6198), .A2(n6478), .ZN(n6490) );
  NAND2_X1 U6015 ( .A1(n6479), .A2(n6477), .ZN(n6198) );
  NAND2_X1 U6016 ( .A1(n6196), .A2(n6197), .ZN(n6477) );
  NAND4_X1 U6017 ( .A1(n6195), .A2(n6194), .A3(n6193), .A4(n6192), .ZN(n6196)
         );
  NAND2_X1 U6018 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[32] ), .A2(n5189), .ZN(
        n6192) );
  NAND2_X1 U6019 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[32] ), .A2(n5154), 
        .ZN(n6193) );
  NAND2_X1 U6020 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[33] ), .A2(n3945), .ZN(
        n6194) );
  AOI21_X1 U6021 ( .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[33] ), .B2(n3946), 
        .A(n6191), .ZN(n6195) );
  NOR2_X1 U6022 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[33] ), .ZN(n6191) );
  NOR2_X1 U6023 ( .A1(n6313), .A2(n6312), .ZN(n6479) );
  NAND4_X1 U6024 ( .A1(n6190), .A2(n6189), .A3(n6188), .A4(n6187), .ZN(n6313)
         );
  NAND2_X1 U6025 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[31] ), .A2(n6298), .ZN(
        n6187) );
  NAND2_X1 U6026 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[31] ), .A2(n5154), 
        .ZN(n6188) );
  NAND2_X1 U6027 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[32] ), .A2(n3945), .ZN(
        n6189) );
  AOI21_X1 U6028 ( .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[32] ), .B2(n3946), 
        .A(n6186), .ZN(n6190) );
  NOR2_X1 U6029 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[32] ), .ZN(n6186) );
  NAND2_X1 U6030 ( .A1(n6216), .A2(n6215), .ZN(n6526) );
  NAND4_X1 U6031 ( .A1(n6209), .A2(n6208), .A3(n6207), .A4(n6206), .ZN(n6216)
         );
  NAND2_X1 U6032 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[38] ), .A2(n3946), 
        .ZN(n6206) );
  NAND2_X1 U6033 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[38] ), .A2(n3945), .ZN(
        n6207) );
  NAND2_X1 U6034 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[37] ), .A2(n6298), .ZN(
        n6208) );
  AOI21_X1 U6035 ( .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[37] ), .B2(n5154), 
        .A(n6205), .ZN(n6209) );
  NOR2_X1 U6036 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[38] ), .ZN(n6205) );
  NAND2_X1 U6037 ( .A1(n6217), .A2(n6218), .ZN(n6518) );
  NAND2_X1 U6038 ( .A1(n6866), .A2(n6865), .ZN(n2940) );
  NAND2_X1 U6039 ( .A1(n7056), .A2(n6864), .ZN(n6865) );
  INV_X1 U6040 ( .A(n6868), .ZN(n6864) );
  NAND2_X1 U6041 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[6] ), .ZN(n6866) );
  NAND2_X1 U6042 ( .A1(n6860), .A2(n6859), .ZN(n2939) );
  NAND2_X1 U6043 ( .A1(n5200), .A2(n6858), .ZN(n6859) );
  INV_X1 U6044 ( .A(n6862), .ZN(n6858) );
  NAND2_X1 U6045 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[7] ), .ZN(n6860) );
  NAND2_X1 U6046 ( .A1(n6991), .A2(rs_id[0]), .ZN(n6985) );
  NAND2_X1 U6047 ( .A1(n6991), .A2(rt_id[3]), .ZN(n6989) );
  NAND2_X1 U6048 ( .A1(n6991), .A2(rt_id[4]), .ZN(n6987) );
  NAND2_X1 U6049 ( .A1(n7005), .A2(n6980), .ZN(n6993) );
  INV_X1 U6050 ( .A(n7060), .ZN(n7005) );
  NAND2_X1 U6051 ( .A1(n6991), .A2(rt_id[2]), .ZN(n6992) );
  AND2_X1 U6052 ( .A1(n5338), .A2(n4354), .ZN(n4872) );
  INV_X1 U6053 ( .A(n4843), .ZN(n4943) );
  OAI211_X1 U6054 ( .C1(n5215), .C2(n6934), .A(n6933), .B(n6932), .ZN(n2725)
         );
  NAND2_X1 U6055 ( .A1(n4107), .A2(n4384), .ZN(n6932) );
  NAND2_X1 U6056 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[31] ), .ZN(n6933) );
  INV_X1 U6057 ( .A(\dp/ids/rp2[31] ), .ZN(n6934) );
  OAI211_X1 U6058 ( .C1(n5215), .C2(n7045), .A(n7044), .B(n7043), .ZN(n2752)
         );
  NAND2_X1 U6059 ( .A1(n5217), .A2(n4412), .ZN(n7043) );
  NAND2_X1 U6060 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[4] ), .ZN(n7044) );
  OAI211_X1 U6061 ( .C1(n5215), .C2(n7050), .A(n7049), .B(n7048), .ZN(n2753)
         );
  NAND2_X1 U6062 ( .A1(n4107), .A2(n4413), .ZN(n7048) );
  NAND2_X1 U6063 ( .A1(n7100), .A2(\dp/op_b_id_ex_int[3] ), .ZN(n7049) );
  OAI211_X1 U6064 ( .C1(n5215), .C2(n6967), .A(n6966), .B(n6965), .ZN(n2726)
         );
  NAND2_X1 U6065 ( .A1(n5216), .A2(n4408), .ZN(n6965) );
  NAND2_X1 U6066 ( .A1(n7100), .A2(\dp/op_b_id_ex_int[30] ), .ZN(n6966) );
  INV_X1 U6067 ( .A(\dp/ids/rp2[30] ), .ZN(n6967) );
  OAI211_X1 U6068 ( .C1(n5215), .C2(n7103), .A(n7102), .B(n7101), .ZN(n2754)
         );
  NAND2_X1 U6069 ( .A1(n5217), .A2(n4414), .ZN(n7101) );
  NAND2_X1 U6070 ( .A1(n7100), .A2(\dp/op_b_id_ex_int[2] ), .ZN(n7102) );
  OAI211_X1 U6071 ( .C1(n6947), .C2(n4362), .A(n6944), .B(n6943), .ZN(n2705)
         );
  NAND2_X1 U6072 ( .A1(n5214), .A2(\dp/ids/rp2[12] ), .ZN(n6943) );
  AOI22_X1 U6073 ( .A1(n3896), .A2(n4392), .B1(n3956), .B2(n4146), .ZN(n6944)
         );
  NAND2_X1 U6074 ( .A1(n5616), .A2(n5613), .ZN(\ctrl_u/n540 ) );
  INV_X1 U6075 ( .A(n5611), .ZN(n5612) );
  OAI211_X1 U6076 ( .C1(n6947), .C2(n4361), .A(n6906), .B(n6905), .ZN(n2706)
         );
  NAND2_X1 U6077 ( .A1(n5214), .A2(\dp/ids/rp2[11] ), .ZN(n6905) );
  AOI22_X1 U6078 ( .A1(n3896), .A2(n4143), .B1(n3956), .B2(n4390), .ZN(n6906)
         );
  NAND2_X1 U6079 ( .A1(n5616), .A2(n5615), .ZN(\ctrl_u/n541 ) );
  NAND2_X1 U6080 ( .A1(n5611), .A2(n5597), .ZN(n5614) );
  INV_X1 U6081 ( .A(n5596), .ZN(n5597) );
  NAND2_X1 U6082 ( .A1(n5610), .A2(n5652), .ZN(n5616) );
  OR4_X1 U6083 ( .A1(n5619), .A2(n5637), .A3(n5609), .A4(n5608), .ZN(n5610) );
  AOI21_X1 U6084 ( .B1(n5607), .B2(n5606), .A(n5605), .ZN(n5609) );
  INV_X1 U6085 ( .A(n5502), .ZN(n5605) );
  INV_X1 U6086 ( .A(n5604), .ZN(n5606) );
  NOR2_X1 U6087 ( .A1(instr_if[30]), .A2(n5560), .ZN(n5649) );
  OAI211_X1 U6088 ( .C1(\intadd_2/SUM[27] ), .C2(n3937), .A(n6408), .B(n6407), 
        .ZN(n2529) );
  OAI211_X1 U6089 ( .C1(\intadd_1/SUM[29] ), .C2(n7066), .A(n6128), .B(n6127), 
        .ZN(n6129) );
  NAND2_X1 U6090 ( .A1(\dp/exs/alu_unit/shifter_out[30] ), .A2(n7083), .ZN(
        n6127) );
  NAND2_X1 U6091 ( .A1(n5108), .A2(n3952), .ZN(n6125) );
  INV_X1 U6092 ( .A(n6124), .ZN(n5108) );
  AOI21_X1 U6093 ( .B1(n6118), .B2(n6141), .A(n6117), .ZN(n6115) );
  INV_X1 U6094 ( .A(n6118), .ZN(n6133) );
  INV_X1 U6095 ( .A(n6117), .ZN(n6123) );
  XNOR2_X1 U6096 ( .A(n6139), .B(n6140), .ZN(n6117) );
  NOR2_X1 U6097 ( .A1(n4962), .A2(n4870), .ZN(n6408) );
  NOR2_X1 U6098 ( .A1(n3873), .A2(n4519), .ZN(n4870) );
  NAND2_X1 U6099 ( .A1(n3928), .A2(\dp/pc_plus4_out_if_int[28] ), .ZN(n6406)
         );
  XNOR2_X1 U6100 ( .A(\intadd_2/n2 ), .B(n5014), .ZN(\intadd_2/SUM[27] ) );
  XNOR2_X1 U6101 ( .A(n4519), .B(n4367), .ZN(n5014) );
  NAND2_X1 U6102 ( .A1(n4056), .A2(n6723), .ZN(n2915) );
  NAND2_X1 U6103 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[31] ), .ZN(n6723) );
  NAND2_X1 U6104 ( .A1(n6756), .A2(n6750), .ZN(n2888) );
  NAND2_X1 U6105 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[58] ), .ZN(n6750) );
  NAND2_X1 U6106 ( .A1(n4057), .A2(n6751), .ZN(n2887) );
  NAND2_X1 U6107 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[59] ), .ZN(n6751) );
  NAND2_X1 U6108 ( .A1(n4057), .A2(n6753), .ZN(n2885) );
  NAND2_X1 U6109 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[61] ), .ZN(n6753) );
  NAND2_X1 U6110 ( .A1(n4056), .A2(n6725), .ZN(n2913) );
  NAND2_X1 U6111 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[33] ), .ZN(n6725) );
  NAND2_X1 U6112 ( .A1(n4057), .A2(n6727), .ZN(n2911) );
  NAND2_X1 U6113 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[35] ), .ZN(n6727) );
  NAND2_X1 U6114 ( .A1(n4056), .A2(n6752), .ZN(n2886) );
  NAND2_X1 U6115 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[60] ), .ZN(n6752) );
  NAND2_X1 U6116 ( .A1(n4055), .A2(n6726), .ZN(n2912) );
  NAND2_X1 U6117 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[34] ), .ZN(n6726) );
  AOI21_X1 U6118 ( .B1(\dp/exs/alu_unit/shifter_out[2] ), .B2(n3954), .A(n5820), .ZN(n7106) );
  OAI211_X1 U6119 ( .C1(\intadd_1/SUM[1] ), .C2(n7066), .A(n5819), .B(n5818), 
        .ZN(n5820) );
  NAND2_X1 U6120 ( .A1(n5817), .A2(n7076), .ZN(n5818) );
  XNOR2_X1 U6121 ( .A(n5816), .B(n5815), .ZN(n5817) );
  INV_X1 U6122 ( .A(n5825), .ZN(n7107) );
  OAI21_X1 U6123 ( .B1(\dp/imm_id_exe_int[2] ), .B2(\dp/npc_id_exe_int[2] ), 
        .A(n5095), .ZN(n5825) );
  INV_X1 U6124 ( .A(n3928), .ZN(n7105) );
  AOI22_X1 U6125 ( .A1(n5134), .A2(\dp/imm_id_int[0] ), .B1(n3978), .B2(
        instr_if[0]), .ZN(n1642) );
  AOI22_X1 U6126 ( .A1(n5134), .A2(\ctrl_u/curr_ak_id ), .B1(n3978), .B2(
        btb_addr_known_if), .ZN(\ctrl_u/n170 ) );
  AOI22_X1 U6127 ( .A1(n5134), .A2(\dp/imm_id_int[8] ), .B1(n3978), .B2(
        instr_if[8]), .ZN(n1634) );
  AOI22_X1 U6128 ( .A1(n5134), .A2(\dp/imm_id_int[7] ), .B1(n3978), .B2(
        instr_if[7]), .ZN(n1635) );
  INV_X1 U6129 ( .A(n7180), .ZN(n279) );
  AOI22_X1 U6130 ( .A1(n5133), .A2(rs_id[0]), .B1(n5179), .B2(instr_if[21]), 
        .ZN(n7180) );
  INV_X1 U6131 ( .A(n7187), .ZN(n283) );
  AOI22_X1 U6132 ( .A1(n5133), .A2(rs_id[4]), .B1(n5180), .B2(instr_if[25]), 
        .ZN(n7187) );
  INV_X1 U6133 ( .A(n5623), .ZN(\ctrl_u/n556 ) );
  AOI22_X1 U6134 ( .A1(\ctrl_u/curr_mul_in_prog ), .A2(n5622), .B1(n5621), 
        .B2(n5620), .ZN(n5623) );
  INV_X1 U6135 ( .A(n7183), .ZN(n282) );
  AOI22_X1 U6136 ( .A1(n5133), .A2(rs_id[3]), .B1(n5180), .B2(instr_if[24]), 
        .ZN(n7183) );
  OAI211_X1 U6137 ( .C1(n6947), .C2(n4376), .A(n6938), .B(n6937), .ZN(n2711)
         );
  NAND2_X1 U6138 ( .A1(n5213), .A2(\dp/ids/rp2[6] ), .ZN(n6937) );
  AOI22_X1 U6139 ( .A1(n3897), .A2(n4141), .B1(n3947), .B2(n4391), .ZN(n6938)
         );
  NAND2_X1 U6140 ( .A1(n3955), .A2(\dp/ids/rp2[18] ), .ZN(n4687) );
  AOI22_X1 U6141 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[18] ), .B1(n4107), .B2(
        n4424), .ZN(n6994) );
  NAND2_X1 U6142 ( .A1(n4682), .A2(\dp/ids/rp2[23] ), .ZN(n4689) );
  AOI22_X1 U6143 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[23] ), .B1(n5217), .B2(
        n4420), .ZN(n6983) );
  NAND2_X1 U6144 ( .A1(n4682), .A2(\dp/ids/rp2[22] ), .ZN(n4693) );
  AOI22_X1 U6145 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[22] ), .B1(n5217), .B2(
        n4443), .ZN(n6984) );
  NAND2_X1 U6146 ( .A1(n4682), .A2(\dp/ids/rp2[19] ), .ZN(n4694) );
  AOI22_X1 U6147 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[19] ), .B1(n5216), .B2(
        n4423), .ZN(n6990) );
  NAND2_X1 U6148 ( .A1(n4682), .A2(\dp/ids/rp2[21] ), .ZN(n4686) );
  AOI22_X1 U6149 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[21] ), .B1(n5217), .B2(
        n4421), .ZN(n6986) );
  NAND2_X1 U6150 ( .A1(n4682), .A2(\dp/ids/rp2[24] ), .ZN(n4685) );
  AOI22_X1 U6151 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[24] ), .B1(n5216), .B2(
        n4419), .ZN(n6982) );
  NAND2_X1 U6152 ( .A1(n3955), .A2(\dp/ids/rp2[20] ), .ZN(n4690) );
  AOI22_X1 U6153 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[20] ), .B1(n4107), .B2(
        n4422), .ZN(n6988) );
  NAND2_X1 U6154 ( .A1(n4682), .A2(\dp/ids/rp2[28] ), .ZN(n4684) );
  AOI22_X1 U6155 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[28] ), .B1(n5216), .B2(
        n4416), .ZN(n6971) );
  NAND2_X1 U6156 ( .A1(n3955), .A2(\dp/ids/rp2[14] ), .ZN(n4695) );
  AOI22_X1 U6157 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[14] ), .B1(n5217), .B2(
        n4426), .ZN(n7011) );
  NAND2_X1 U6158 ( .A1(n3955), .A2(\dp/ids/rp2[26] ), .ZN(n4692) );
  AOI22_X1 U6159 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[26] ), .B1(n5216), .B2(
        n4418), .ZN(n6977) );
  NAND2_X1 U6160 ( .A1(n4682), .A2(\dp/ids/rp2[29] ), .ZN(n4691) );
  AOI22_X1 U6161 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[29] ), .B1(n4107), .B2(
        n4415), .ZN(n6969) );
  NAND2_X1 U6162 ( .A1(n3955), .A2(\dp/ids/rp2[27] ), .ZN(n4688) );
  AOI22_X1 U6163 ( .A1(n5128), .A2(\dp/op_b_id_ex_int[27] ), .B1(n4107), .B2(
        n4417), .ZN(n6973) );
  OAI21_X1 U6164 ( .B1(n3934), .B2(n5487), .A(n5486), .ZN(\ctrl_u/n507 ) );
  OAI21_X1 U6165 ( .B1(n3934), .B2(n5485), .A(n5484), .ZN(\ctrl_u/n506 ) );
  NOR2_X1 U6166 ( .A1(n5483), .A2(n5482), .ZN(n5579) );
  NAND4_X1 U6167 ( .A1(n7293), .A2(instr_if[4]), .A3(n5530), .A4(n7277), .ZN(
        n5482) );
  OAI21_X1 U6168 ( .B1(\ctrl_u/curr_id[25] ), .B2(n5652), .A(n5642), .ZN(
        \ctrl_u/n335 ) );
  OAI21_X1 U6169 ( .B1(n5467), .B2(n5438), .A(n5499), .ZN(n5639) );
  OAI21_X1 U6170 ( .B1(n7284), .B2(n7278), .A(n5437), .ZN(n5438) );
  AOI21_X1 U6171 ( .B1(instr_if[0]), .B2(n7284), .A(n5596), .ZN(n5437) );
  NAND2_X1 U6172 ( .A1(instr_if[5]), .A2(n5585), .ZN(n5467) );
  AOI211_X1 U6173 ( .C1(n5638), .C2(instr_if[16]), .A(n5637), .B(n5636), .ZN(
        n5640) );
  NAND4_X1 U6174 ( .A1(n5635), .A2(n5634), .A3(n5633), .A4(n5632), .ZN(n5636)
         );
  OAI21_X1 U6175 ( .B1(instr_if[27]), .B2(n5631), .A(instr_if[26]), .ZN(n5632)
         );
  INV_X1 U6176 ( .A(n5630), .ZN(n5631) );
  NOR2_X1 U6177 ( .A1(n5629), .A2(n5628), .ZN(n5634) );
  NOR3_X1 U6178 ( .A1(instr_if[28]), .A2(instr_if[29]), .A3(n5627), .ZN(n5628)
         );
  AOI22_X1 U6179 ( .A1(n5647), .A2(instr_if[28]), .B1(n5590), .B2(n5587), .ZN(
        n5635) );
  OAI21_X1 U6180 ( .B1(\ctrl_u/curr_id[6] ), .B2(n5652), .A(n5603), .ZN(
        \ctrl_u/n402 ) );
  NOR4_X1 U6181 ( .A1(n5637), .A2(n5600), .A3(n5611), .A4(n7296), .ZN(n5601)
         );
  NOR2_X1 U6182 ( .A1(n5595), .A2(n5594), .ZN(n5611) );
  NOR3_X1 U6183 ( .A1(n5608), .A2(n5593), .A3(n5592), .ZN(n5602) );
  OAI21_X1 U6184 ( .B1(n5591), .B2(n5590), .A(n5630), .ZN(n5592) );
  AOI21_X1 U6185 ( .B1(instr_if[31]), .B2(n5589), .A(n5607), .ZN(n5593) );
  AOI21_X1 U6186 ( .B1(instr_if[27]), .B2(n5588), .A(n5587), .ZN(n5607) );
  INV_X1 U6187 ( .A(n5445), .ZN(n5587) );
  NOR2_X1 U6188 ( .A1(instr_if[28]), .A2(n5560), .ZN(n5588) );
  NOR2_X1 U6189 ( .A1(n5586), .A2(n5594), .ZN(n5608) );
  AND3_X1 U6190 ( .A1(n7287), .A2(n5585), .A3(n7281), .ZN(n5586) );
  NOR2_X1 U6191 ( .A1(n5497), .A2(n7279), .ZN(n5585) );
  OAI211_X1 U6192 ( .C1(n6947), .C2(n4364), .A(n6946), .B(n6945), .ZN(n2703)
         );
  NAND2_X1 U6193 ( .A1(n5213), .A2(\dp/ids/rp2[14] ), .ZN(n6945) );
  AOI22_X1 U6194 ( .A1(n3898), .A2(n4146), .B1(n5211), .B2(n4395), .ZN(n6946)
         );
  OAI211_X1 U6195 ( .C1(n6947), .C2(n4375), .A(n6902), .B(n6901), .ZN(n2710)
         );
  NAND2_X1 U6196 ( .A1(n5214), .A2(\dp/ids/rp2[7] ), .ZN(n6901) );
  AOI22_X1 U6197 ( .A1(n3897), .A2(n4142), .B1(n5211), .B2(n4389), .ZN(n6902)
         );
  OAI211_X1 U6198 ( .C1(n6947), .C2(n4363), .A(n6908), .B(n6907), .ZN(n2704)
         );
  NAND2_X1 U6199 ( .A1(n5213), .A2(\dp/ids/rp2[13] ), .ZN(n6907) );
  AOI22_X1 U6200 ( .A1(n3898), .A2(n4390), .B1(n5211), .B2(n4144), .ZN(n6908)
         );
  OAI211_X1 U6201 ( .C1(n6947), .C2(n4374), .A(n6940), .B(n6939), .ZN(n2709)
         );
  NAND2_X1 U6202 ( .A1(n5214), .A2(\dp/ids/rp2[8] ), .ZN(n6939) );
  AOI22_X1 U6203 ( .A1(n3896), .A2(n4391), .B1(n5211), .B2(n4145), .ZN(n6940)
         );
  OAI22_X1 U6204 ( .A1(n7058), .A2(n6894), .B1(n4049), .B2(n613), .ZN(n2978)
         );
  OAI22_X1 U6205 ( .A1(n4051), .A2(n644), .B1(n7058), .B2(n6758), .ZN(n2947)
         );
  INV_X1 U6206 ( .A(n6722), .ZN(n6758) );
  OAI22_X1 U6207 ( .A1(n4049), .A2(n4262), .B1(n4047), .B2(n7052), .ZN(n2719)
         );
  AOI21_X1 U6208 ( .B1(\dp/imm_id_int[2] ), .B2(n4357), .A(n6935), .ZN(n7052)
         );
  NOR2_X1 U6209 ( .A1(n7103), .A2(n4357), .ZN(n6935) );
  AOI21_X1 U6210 ( .B1(instr_if[0]), .B2(n5480), .A(n5550), .ZN(n5428) );
  NOR3_X1 U6211 ( .A1(n5490), .A2(n5548), .A3(n3962), .ZN(n5550) );
  INV_X1 U6212 ( .A(n7284), .ZN(n5595) );
  OAI22_X1 U6213 ( .A1(n4050), .A2(n4263), .B1(n4048), .B2(n7054), .ZN(n2720)
         );
  AOI21_X1 U6214 ( .B1(\dp/ids/rp2[1] ), .B2(b_selector_id), .A(n6895), .ZN(
        n7054) );
  NOR2_X1 U6215 ( .A1(n4476), .A2(b_selector_id), .ZN(n6895) );
  OAI21_X1 U6216 ( .B1(n5182), .B2(n5555), .A(n5554), .ZN(\ctrl_u/n544 ) );
  NAND2_X1 U6217 ( .A1(n4057), .A2(n6748), .ZN(n2890) );
  NAND2_X1 U6218 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[56] ), .ZN(n6748) );
  OAI211_X1 U6219 ( .C1(n6947), .C2(n4373), .A(n6904), .B(n6903), .ZN(n2708)
         );
  NAND2_X1 U6220 ( .A1(n5213), .A2(\dp/ids/rp2[9] ), .ZN(n6903) );
  AOI22_X1 U6221 ( .A1(n3896), .A2(n4389), .B1(n3947), .B2(n4143), .ZN(n6904)
         );
  OAI211_X1 U6222 ( .C1(n6947), .C2(n4372), .A(n6942), .B(n6941), .ZN(n2707)
         );
  NAND2_X1 U6223 ( .A1(n5213), .A2(\dp/ids/rp2[10] ), .ZN(n6941) );
  AOI22_X1 U6224 ( .A1(n3898), .A2(n4145), .B1(n3947), .B2(n4392), .ZN(n6942)
         );
  OAI211_X1 U6225 ( .C1(n6947), .C2(n4368), .A(n6910), .B(n6909), .ZN(n2702)
         );
  NAND2_X1 U6226 ( .A1(n5214), .A2(\dp/ids/rp2[15] ), .ZN(n6909) );
  AOI22_X1 U6227 ( .A1(n3897), .A2(n4144), .B1(n3947), .B2(n4394), .ZN(n6910)
         );
  OAI22_X1 U6228 ( .A1(n4047), .A2(n6838), .B1(n4050), .B2(n629), .ZN(n2962)
         );
  AOI21_X1 U6229 ( .B1(\dp/ids/rp1[16] ), .B2(n4136), .A(n6836), .ZN(n6838) );
  NOR2_X1 U6230 ( .A1(n4136), .A2(n374), .ZN(n6836) );
  OAI22_X1 U6231 ( .A1(n4047), .A2(n6841), .B1(n4050), .B2(n628), .ZN(n2963)
         );
  AOI21_X1 U6232 ( .B1(\dp/ids/rp1[15] ), .B2(n4136), .A(n6839), .ZN(n6841) );
  NOR2_X1 U6233 ( .A1(n4136), .A2(n373), .ZN(n6839) );
  NOR2_X1 U6234 ( .A1(n5619), .A2(n4772), .ZN(n5344) );
  NAND2_X1 U6235 ( .A1(n4774), .A2(n4773), .ZN(n4772) );
  NAND2_X1 U6236 ( .A1(n3912), .A2(\ctrl_u/curr_mul_end_wb ), .ZN(n4773) );
  INV_X1 U6237 ( .A(n5158), .ZN(n4774) );
  AOI211_X1 U6238 ( .C1(n5647), .C2(n5466), .A(n5629), .B(n5600), .ZN(n5474)
         );
  INV_X1 U6239 ( .A(n5465), .ZN(n5600) );
  NOR2_X1 U6240 ( .A1(n5514), .A2(n5590), .ZN(n5629) );
  INV_X1 U6241 ( .A(n5494), .ZN(n5466) );
  OAI211_X1 U6242 ( .C1(n5462), .C2(n5461), .A(n5460), .B(n5459), .ZN(n5463)
         );
  INV_X1 U6243 ( .A(n7282), .ZN(n5459) );
  OAI21_X1 U6244 ( .B1(instr_if[4]), .B2(instr_if[0]), .A(n5596), .ZN(n5460)
         );
  OAI21_X1 U6245 ( .B1(n7283), .B2(n7279), .A(n7277), .ZN(n5461) );
  NOR3_X1 U6246 ( .A1(instr_if[3]), .A2(instr_if[0]), .A3(n7278), .ZN(n5462)
         );
  OAI21_X1 U6247 ( .B1(n7284), .B2(n7278), .A(n7285), .ZN(n5464) );
  OAI21_X1 U6248 ( .B1(n5027), .B2(\ctrl_u/n555 ), .A(n4867), .ZN(n4876) );
  NAND2_X1 U6249 ( .A1(n7274), .A2(rst_mem_wb_regs), .ZN(n5350) );
  NOR2_X1 U6250 ( .A1(n5347), .A2(n5346), .ZN(n5354) );
  NOR2_X1 U6251 ( .A1(n5339), .A2(n4867), .ZN(n4866) );
  AND2_X1 U6252 ( .A1(n5338), .A2(n4323), .ZN(n4868) );
  INV_X1 U6253 ( .A(n5417), .ZN(n5617) );
  OAI22_X1 U6254 ( .A1(n7058), .A2(n6889), .B1(n4049), .B2(n614), .ZN(n2977)
         );
  NAND2_X1 U6255 ( .A1(n4971), .A2(n4894), .ZN(n4970) );
  NAND2_X1 U6256 ( .A1(n3884), .A2(n4895), .ZN(n4894) );
  AOI21_X1 U6257 ( .B1(n6071), .B2(n7076), .A(n6070), .ZN(n6419) );
  OAI211_X1 U6258 ( .C1(\intadd_1/SUM[24] ), .C2(n7066), .A(n6069), .B(n6068), 
        .ZN(n6070) );
  NAND2_X1 U6259 ( .A1(n5110), .A2(n3952), .ZN(n6066) );
  INV_X1 U6260 ( .A(n6065), .ZN(n5110) );
  NAND2_X1 U6261 ( .A1(\dp/exs/alu_unit/shifter_out[25] ), .A2(n3954), .ZN(
        n6069) );
  XNOR2_X1 U6262 ( .A(n6074), .B(n6073), .ZN(n6064) );
  XNOR2_X1 U6263 ( .A(n4137), .B(n4211), .ZN(n4748) );
  OAI21_X1 U6264 ( .B1(n3957), .B2(n4747), .A(n4746), .ZN(n4749) );
  NAND2_X1 U6265 ( .A1(n4979), .A2(n4898), .ZN(n4978) );
  NAND2_X1 U6266 ( .A1(n3884), .A2(n4899), .ZN(n4898) );
  OAI211_X1 U6267 ( .C1(n7066), .C2(\intadd_1/SUM[27] ), .A(n6109), .B(n6108), 
        .ZN(n6110) );
  NAND2_X1 U6268 ( .A1(\dp/exs/alu_unit/shifter_out[28] ), .A2(n3954), .ZN(
        n6108) );
  NAND2_X1 U6269 ( .A1(n5113), .A2(n3952), .ZN(n6106) );
  INV_X1 U6270 ( .A(n6105), .ZN(n5113) );
  XNOR2_X1 U6271 ( .A(n6136), .B(n6135), .ZN(n6104) );
  AOI22_X1 U6272 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[28] ), .A2(n3945), .B1(
        n6327), .B2(n4286), .ZN(n6101) );
  AOI22_X1 U6273 ( .A1(n3946), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[28] ), 
        .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[27] ), .B2(n6326), .ZN(n6102)
         );
  INV_X1 U6274 ( .A(\dp/exs/alu_unit/mult/a_shiftn[27] ), .ZN(n6103) );
  AOI22_X1 U6275 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[27] ), .A2(n3945), .B1(
        n6327), .B2(n4404), .ZN(n6091) );
  AOI22_X1 U6276 ( .A1(n3946), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[27] ), 
        .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[26] ), .B2(n6326), .ZN(n6092)
         );
  INV_X1 U6277 ( .A(\dp/exs/alu_unit/mult/a_shiftn[26] ), .ZN(n6093) );
  NAND2_X1 U6278 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[26] ), .ZN(n6094)
         );
  AOI22_X1 U6279 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[27] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[27] ), .ZN(n6095) );
  NAND2_X1 U6280 ( .A1(n4896), .A2(n4975), .ZN(n4974) );
  NAND2_X1 U6281 ( .A1(n3884), .A2(n4897), .ZN(n4896) );
  AOI21_X1 U6282 ( .B1(n6086), .B2(n7076), .A(n6085), .ZN(n6418) );
  OAI211_X1 U6283 ( .C1(\intadd_1/SUM[25] ), .C2(n7066), .A(n6084), .B(n6083), 
        .ZN(n6085) );
  NOR2_X1 U6284 ( .A1(n4236), .A2(op_type_exe[1]), .ZN(n5751) );
  NAND2_X1 U6285 ( .A1(\dp/exs/alu_unit/shifter_out[26] ), .A2(n3954), .ZN(
        n6084) );
  OAI21_X1 U6286 ( .B1(n621), .B2(n5175), .A(n7236), .ZN(
        \dp/exs/a_shift_int[8] ) );
  INV_X1 U6287 ( .A(n7235), .ZN(n7236) );
  OAI21_X1 U6288 ( .B1(n619), .B2(n5174), .A(n7240), .ZN(
        \dp/exs/a_shift_int[6] ) );
  INV_X1 U6289 ( .A(n7239), .ZN(n7240) );
  OAI21_X1 U6290 ( .B1(n617), .B2(n3949), .A(n7244), .ZN(
        \dp/exs/a_shift_int[4] ) );
  INV_X1 U6291 ( .A(n7243), .ZN(n7244) );
  OAI21_X1 U6292 ( .B1(n625), .B2(n3949), .A(n7228), .ZN(
        \dp/exs/a_shift_int[12] ) );
  INV_X1 U6293 ( .A(n7227), .ZN(n7228) );
  OAI21_X1 U6294 ( .B1(n631), .B2(n3949), .A(n7216), .ZN(
        \dp/exs/a_shift_int[18] ) );
  INV_X1 U6295 ( .A(n7215), .ZN(n7216) );
  OAI21_X1 U6296 ( .B1(n629), .B2(n5175), .A(n7220), .ZN(
        \dp/exs/a_shift_int[16] ) );
  INV_X1 U6297 ( .A(n7219), .ZN(n7220) );
  OAI21_X1 U6298 ( .B1(n624), .B2(n3949), .A(n7230), .ZN(
        \dp/exs/a_shift_int[11] ) );
  INV_X1 U6299 ( .A(n7229), .ZN(n7230) );
  OAI21_X1 U6300 ( .B1(n628), .B2(n3949), .A(n7222), .ZN(
        \dp/exs/a_shift_int[15] ) );
  INV_X1 U6301 ( .A(n7221), .ZN(n7222) );
  OAI21_X1 U6302 ( .B1(n626), .B2(n3949), .A(n7226), .ZN(
        \dp/exs/a_shift_int[13] ) );
  INV_X1 U6303 ( .A(n7225), .ZN(n7226) );
  OAI21_X1 U6304 ( .B1(n640), .B2(n3949), .A(n7198), .ZN(
        \dp/exs/a_shift_int[27] ) );
  INV_X1 U6305 ( .A(n7197), .ZN(n7198) );
  OAI21_X1 U6306 ( .B1(n636), .B2(n5174), .A(n7206), .ZN(
        \dp/exs/a_shift_int[23] ) );
  INV_X1 U6307 ( .A(n7205), .ZN(n7206) );
  OAI21_X1 U6308 ( .B1(n643), .B2(n5175), .A(n7192), .ZN(
        \dp/exs/a_shift_int[30] ) );
  INV_X1 U6309 ( .A(n7191), .ZN(n7192) );
  OAI21_X1 U6310 ( .B1(n632), .B2(n5175), .A(n7214), .ZN(
        \dp/exs/a_shift_int[19] ) );
  INV_X1 U6311 ( .A(n7213), .ZN(n7214) );
  OAI21_X1 U6312 ( .B1(n613), .B2(n3949), .A(n7252), .ZN(
        \dp/exs/a_shift_int[0] ) );
  INV_X1 U6313 ( .A(n7251), .ZN(n7252) );
  OAI21_X1 U6314 ( .B1(n615), .B2(n5174), .A(n7248), .ZN(
        \dp/exs/a_shift_int[2] ) );
  INV_X1 U6315 ( .A(n7247), .ZN(n7248) );
  OAI21_X1 U6316 ( .B1(n614), .B2(n3949), .A(n7250), .ZN(
        \dp/exs/a_shift_int[1] ) );
  INV_X1 U6317 ( .A(n7249), .ZN(n7250) );
  OAI21_X1 U6318 ( .B1(n622), .B2(n5174), .A(n7234), .ZN(
        \dp/exs/a_shift_int[9] ) );
  INV_X1 U6319 ( .A(n7233), .ZN(n7234) );
  OAI21_X1 U6320 ( .B1(n620), .B2(n3949), .A(n7238), .ZN(
        \dp/exs/a_shift_int[7] ) );
  INV_X1 U6321 ( .A(n7237), .ZN(n7238) );
  OAI21_X1 U6322 ( .B1(n616), .B2(n3949), .A(n7246), .ZN(
        \dp/exs/a_shift_int[3] ) );
  INV_X1 U6323 ( .A(n7245), .ZN(n7246) );
  OAI21_X1 U6324 ( .B1(n642), .B2(n3949), .A(n7194), .ZN(
        \dp/exs/a_shift_int[29] ) );
  INV_X1 U6325 ( .A(n7193), .ZN(n7194) );
  OAI21_X1 U6326 ( .B1(n635), .B2(n5174), .A(n7208), .ZN(
        \dp/exs/a_shift_int[22] ) );
  INV_X1 U6327 ( .A(n7207), .ZN(n7208) );
  OAI21_X1 U6328 ( .B1(n639), .B2(n3949), .A(n7200), .ZN(
        \dp/exs/a_shift_int[26] ) );
  INV_X1 U6329 ( .A(n7199), .ZN(n7200) );
  OAI21_X1 U6330 ( .B1(n634), .B2(n5174), .A(n7210), .ZN(
        \dp/exs/a_shift_int[21] ) );
  INV_X1 U6331 ( .A(n7209), .ZN(n7210) );
  OAI21_X1 U6332 ( .B1(n641), .B2(n3949), .A(n7196), .ZN(
        \dp/exs/a_shift_int[28] ) );
  INV_X1 U6333 ( .A(n7195), .ZN(n7196) );
  OAI21_X1 U6334 ( .B1(n638), .B2(n3949), .A(n7202), .ZN(
        \dp/exs/a_shift_int[25] ) );
  INV_X1 U6335 ( .A(n7201), .ZN(n7202) );
  OAI21_X1 U6336 ( .B1(n627), .B2(n3949), .A(n7224), .ZN(
        \dp/exs/a_shift_int[14] ) );
  INV_X1 U6337 ( .A(n7223), .ZN(n7224) );
  OAI21_X1 U6338 ( .B1(n618), .B2(n5175), .A(n7242), .ZN(
        \dp/exs/a_shift_int[5] ) );
  INV_X1 U6339 ( .A(n7241), .ZN(n7242) );
  OAI21_X1 U6340 ( .B1(n623), .B2(n5175), .A(n7232), .ZN(
        \dp/exs/a_shift_int[10] ) );
  INV_X1 U6341 ( .A(n7231), .ZN(n7232) );
  OAI21_X1 U6342 ( .B1(n630), .B2(n5175), .A(n7218), .ZN(
        \dp/exs/a_shift_int[17] ) );
  INV_X1 U6343 ( .A(n7217), .ZN(n7218) );
  OAI21_X1 U6344 ( .B1(n7260), .B2(n4260), .A(n7255), .ZN(n110) );
  INV_X1 U6345 ( .A(n7254), .ZN(n7255) );
  OAI21_X1 U6346 ( .B1(n7260), .B2(n4261), .A(n7256), .ZN(n103) );
  OAI21_X1 U6347 ( .B1(n644), .B2(n5174), .A(n7190), .ZN(
        \dp/exs/a_shift_int[31] ) );
  INV_X1 U6348 ( .A(n7189), .ZN(n7190) );
  OAI21_X1 U6349 ( .B1(n637), .B2(n5175), .A(n7204), .ZN(
        \dp/exs/a_shift_int[24] ) );
  INV_X1 U6350 ( .A(n7203), .ZN(n7204) );
  OAI21_X1 U6351 ( .B1(n633), .B2(n5174), .A(n7212), .ZN(
        \dp/exs/a_shift_int[20] ) );
  INV_X1 U6352 ( .A(n7211), .ZN(n7212) );
  XNOR2_X1 U6353 ( .A(n6089), .B(n6090), .ZN(n6081) );
  OAI211_X1 U6354 ( .C1(n3930), .C2(n4065), .A(n6080), .B(n6079), .ZN(n6090)
         );
  NAND2_X1 U6355 ( .A1(n3943), .A2(\dp/a_neg_mult_id_exe_int[25] ), .ZN(n6079)
         );
  AOI22_X1 U6356 ( .A1(\dp/a_neg_mult_id_exe_int[26] ), .A2(n3939), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[26] ), .ZN(n6080) );
  OAI211_X1 U6357 ( .C1(n6078), .C2(n6328), .A(n6077), .B(n6076), .ZN(n6089)
         );
  AOI22_X1 U6358 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[26] ), .A2(n3945), .B1(
        n6327), .B2(n4274), .ZN(n6076) );
  AOI22_X1 U6359 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[25] ), .A2(n6326), 
        .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[26] ), .B2(n3946), .ZN(n6077)
         );
  INV_X1 U6360 ( .A(\dp/exs/alu_unit/mult/a_shiftn[25] ), .ZN(n6078) );
  OAI211_X1 U6361 ( .C1(n3930), .C2(n4062), .A(n6063), .B(n6062), .ZN(n6073)
         );
  NAND2_X1 U6362 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[24] ), .ZN(n6062)
         );
  AOI22_X1 U6363 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[25] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[25] ), .ZN(n6063) );
  OAI211_X1 U6364 ( .C1(n6061), .C2(n6060), .A(n6059), .B(n6058), .ZN(n6074)
         );
  AOI22_X1 U6365 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[24] ), .A2(n5189), .B1(
        n6327), .B2(n4273), .ZN(n6058) );
  AOI22_X1 U6366 ( .A1(n3945), .A2(\dp/exs/alu_unit/mult/a_shiftn[25] ), .B1(
        \dp/exs/alu_unit/mult/neg_a_shiftn[24] ), .B2(n5154), .ZN(n6059) );
  INV_X1 U6367 ( .A(\dp/exs/alu_unit/mult/neg_a_shiftn[25] ), .ZN(n6060) );
  NOR2_X1 U6368 ( .A1(n4861), .A2(n4860), .ZN(n4859) );
  INV_X1 U6369 ( .A(n5028), .ZN(n4860) );
  AOI22_X1 U6370 ( .A1(n5030), .A2(n5032), .B1(n5033), .B2(n5036), .ZN(n5028)
         );
  NAND2_X1 U6371 ( .A1(n5064), .A2(n5037), .ZN(n5036) );
  INV_X1 U6372 ( .A(n6040), .ZN(n5037) );
  NOR2_X1 U6373 ( .A1(n5029), .A2(n4858), .ZN(n4857) );
  INV_X1 U6374 ( .A(n4863), .ZN(n4858) );
  NAND2_X1 U6375 ( .A1(n4902), .A2(n4864), .ZN(n4863) );
  INV_X1 U6376 ( .A(n4904), .ZN(n4864) );
  AOI21_X1 U6377 ( .B1(n4905), .B2(n5006), .A(n4324), .ZN(n4904) );
  OAI211_X1 U6378 ( .C1(n3930), .C2(n4076), .A(n5990), .B(n5989), .ZN(n6005)
         );
  NAND2_X1 U6379 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[19] ), .ZN(n5989)
         );
  AOI22_X1 U6380 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[20] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[20] ), .ZN(n5990) );
  OAI211_X1 U6381 ( .C1(n6328), .C2(n5993), .A(n5992), .B(n5991), .ZN(n6004)
         );
  AOI22_X1 U6382 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[20] ), .A2(n3946), 
        .B1(n6327), .B2(n4269), .ZN(n5991) );
  AOI22_X1 U6383 ( .A1(n3945), .A2(\dp/exs/alu_unit/mult/a_shiftn[20] ), .B1(
        \dp/exs/alu_unit/mult/neg_a_shiftn[19] ), .B2(n6326), .ZN(n5992) );
  INV_X1 U6384 ( .A(\dp/exs/alu_unit/mult/a_shiftn[19] ), .ZN(n5993) );
  NAND2_X1 U6385 ( .A1(n5987), .A2(n5986), .ZN(n5006) );
  INV_X1 U6386 ( .A(n5007), .ZN(n4905) );
  OR2_X1 U6387 ( .A1(n5987), .A2(n5986), .ZN(n5007) );
  OAI211_X1 U6388 ( .C1(n3930), .C2(n4075), .A(n5973), .B(n5972), .ZN(n5986)
         );
  NAND2_X1 U6389 ( .A1(n3943), .A2(\dp/a_neg_mult_id_exe_int[18] ), .ZN(n5972)
         );
  AOI22_X1 U6390 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[19] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[19] ), .ZN(n5973) );
  OAI211_X1 U6391 ( .C1(n6061), .C2(n5976), .A(n5975), .B(n5974), .ZN(n5987)
         );
  AOI22_X1 U6392 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[18] ), .A2(n5189), .B1(
        n6327), .B2(n4268), .ZN(n5974) );
  AOI22_X1 U6393 ( .A1(n3945), .A2(\dp/exs/alu_unit/mult/a_shiftn[19] ), .B1(
        \dp/exs/alu_unit/mult/neg_a_shiftn[18] ), .B2(n6326), .ZN(n5975) );
  INV_X1 U6394 ( .A(\dp/exs/alu_unit/mult/neg_a_shiftn[19] ), .ZN(n5976) );
  NOR2_X1 U6395 ( .A1(n5030), .A2(n5033), .ZN(n5029) );
  AOI21_X1 U6396 ( .B1(n5035), .B2(n5064), .A(n5034), .ZN(n5033) );
  INV_X1 U6397 ( .A(n6039), .ZN(n5034) );
  OAI211_X1 U6398 ( .C1(n3930), .C2(n4078), .A(n6035), .B(n6034), .ZN(n6039)
         );
  NAND2_X1 U6399 ( .A1(n3943), .A2(\dp/a_neg_mult_id_exe_int[22] ), .ZN(n6034)
         );
  AOI22_X1 U6400 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[23] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[23] ), .ZN(n6035) );
  NOR2_X1 U6401 ( .A1(n4206), .A2(n6040), .ZN(n5035) );
  INV_X1 U6402 ( .A(n5031), .ZN(n5030) );
  OAI21_X1 U6403 ( .B1(n5032), .B2(n4206), .A(n6040), .ZN(n5031) );
  OAI211_X1 U6404 ( .C1(n6061), .C2(n6033), .A(n6032), .B(n6031), .ZN(n6040)
         );
  AOI22_X1 U6405 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[22] ), .A2(n5189), .B1(
        n6327), .B2(n4272), .ZN(n6031) );
  AOI22_X1 U6406 ( .A1(n3945), .A2(\dp/exs/alu_unit/mult/a_shiftn[23] ), .B1(
        \dp/exs/alu_unit/mult/neg_a_shiftn[22] ), .B2(n5154), .ZN(n6032) );
  INV_X1 U6407 ( .A(\dp/exs/alu_unit/mult/neg_a_shiftn[23] ), .ZN(n6033) );
  INV_X1 U6408 ( .A(n5188), .ZN(n6061) );
  NOR2_X1 U6409 ( .A1(n6021), .A2(n6020), .ZN(n5068) );
  AND2_X1 U6410 ( .A1(n6029), .A2(n6030), .ZN(n5066) );
  OAI211_X1 U6411 ( .C1(n3930), .C2(n4077), .A(n6024), .B(n6023), .ZN(n6030)
         );
  NAND2_X1 U6412 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[21] ), .ZN(n6023)
         );
  AOI22_X1 U6413 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[22] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[22] ), .ZN(n6024) );
  AOI22_X1 U6414 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[22] ), .A2(n3945), .B1(
        n6327), .B2(n4271), .ZN(n6025) );
  AOI22_X1 U6415 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[21] ), .A2(n6298), .B1(
        \dp/exs/alu_unit/mult/neg_a_shiftn[22] ), .B2(n3946), .ZN(n6026) );
  INV_X1 U6416 ( .A(n5067), .ZN(n5065) );
  NAND2_X1 U6417 ( .A1(n6021), .A2(n6020), .ZN(n5067) );
  OAI211_X1 U6418 ( .C1(n3930), .C2(n4086), .A(n6007), .B(n6006), .ZN(n6020)
         );
  NAND2_X1 U6419 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[20] ), .ZN(n6006)
         );
  AOI22_X1 U6420 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[21] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[21] ), .ZN(n6007) );
  OAI211_X1 U6421 ( .C1(n6328), .C2(n6010), .A(n6009), .B(n6008), .ZN(n6021)
         );
  AOI22_X1 U6422 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[21] ), .A2(n3945), .B1(
        n6327), .B2(n4270), .ZN(n6008) );
  AOI22_X1 U6423 ( .A1(n3946), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[21] ), 
        .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[20] ), .B2(n6326), .ZN(n6009)
         );
  INV_X1 U6424 ( .A(\dp/exs/alu_unit/mult/a_shiftn[20] ), .ZN(n6010) );
  NAND2_X1 U6425 ( .A1(n5970), .A2(n5971), .ZN(n4800) );
  NAND2_X1 U6426 ( .A1(n5969), .A2(n4310), .ZN(n4801) );
  OAI211_X1 U6427 ( .C1(n3930), .C2(n4085), .A(n5959), .B(n5958), .ZN(n5971)
         );
  NAND2_X1 U6428 ( .A1(n3919), .A2(\dp/a_neg_mult_id_exe_int[17] ), .ZN(n5958)
         );
  AOI22_X1 U6429 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[18] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[18] ), .ZN(n5959) );
  NOR2_X1 U6430 ( .A1(n4786), .A2(n4814), .ZN(n4785) );
  INV_X1 U6431 ( .A(n5102), .ZN(n5101) );
  OAI21_X1 U6432 ( .B1(n5103), .B2(n4106), .A(n5956), .ZN(n5102) );
  INV_X1 U6433 ( .A(n5107), .ZN(n5103) );
  AOI21_X1 U6434 ( .B1(n5106), .B2(n5107), .A(n5105), .ZN(n5104) );
  INV_X1 U6435 ( .A(n5955), .ZN(n5105) );
  NOR2_X1 U6436 ( .A1(n5757), .A2(n5756), .ZN(n5107) );
  NOR2_X1 U6437 ( .A1(n4106), .A2(n5956), .ZN(n5106) );
  NAND4_X1 U6438 ( .A1(n5750), .A2(n5749), .A3(n5748), .A4(n5747), .ZN(n5757)
         );
  NAND2_X1 U6439 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[15] ), .A2(n6298), .ZN(
        n5747) );
  NAND2_X1 U6440 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[16] ), .A2(n5188), 
        .ZN(n5748) );
  NAND2_X1 U6441 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[16] ), .A2(n3945), .ZN(
        n5749) );
  AOI21_X1 U6442 ( .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[15] ), .B2(n5154), 
        .A(n5746), .ZN(n5750) );
  NOR2_X1 U6443 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[16] ), .ZN(n5746) );
  NAND2_X1 U6444 ( .A1(n4950), .A2(n4951), .ZN(n4763) );
  AOI22_X1 U6445 ( .A1(n4955), .A2(n4957), .B1(n4952), .B2(n4954), .ZN(n4951)
         );
  INV_X1 U6446 ( .A(n4990), .ZN(n4954) );
  AOI21_X1 U6447 ( .B1(n4953), .B2(n4990), .A(n4958), .ZN(n4952) );
  INV_X1 U6448 ( .A(n4991), .ZN(n4953) );
  INV_X1 U6449 ( .A(n4956), .ZN(n4955) );
  OAI21_X1 U6450 ( .B1(n4957), .B2(n4991), .A(n5939), .ZN(n4956) );
  NAND2_X1 U6451 ( .A1(n4990), .A2(n4958), .ZN(n4957) );
  NAND4_X1 U6452 ( .A1(n5745), .A2(n5744), .A3(n5743), .A4(n5742), .ZN(n5940)
         );
  NAND2_X1 U6453 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[13] ), .A2(n5189), .ZN(
        n5742) );
  NAND2_X1 U6454 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[13] ), .A2(n6326), 
        .ZN(n5743) );
  NAND2_X1 U6455 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[14] ), .A2(n3946), 
        .ZN(n5744) );
  AOI21_X1 U6456 ( .B1(\dp/exs/alu_unit/mult/a_shiftn[14] ), .B2(n3945), .A(
        n5741), .ZN(n5745) );
  NOR2_X1 U6457 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[14] ), .ZN(n5741) );
  NOR2_X1 U6458 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[13] ), .ZN(n5688) );
  INV_X1 U6459 ( .A(n5886), .ZN(n5734) );
  INV_X1 U6460 ( .A(n5885), .ZN(n5729) );
  NAND2_X1 U6461 ( .A1(n5185), .A2(\dp/a_mult_id_exe_int[7] ), .ZN(n5727) );
  NAND2_X1 U6462 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[7] ), .ZN(n5728)
         );
  INV_X1 U6463 ( .A(n5719), .ZN(n5854) );
  NOR2_X1 U6464 ( .A1(n3900), .A2(\dp/a_mult_id_exe_int[1] ), .ZN(n6468) );
  AOI21_X1 U6465 ( .B1(n5153), .B2(n5715), .A(n5714), .ZN(n5717) );
  NOR2_X1 U6466 ( .A1(n3900), .A2(\dp/a_mult_id_exe_int[0] ), .ZN(n5714) );
  AOI21_X1 U6467 ( .B1(n593), .B2(n4230), .A(n5713), .ZN(n5715) );
  OAI21_X1 U6468 ( .B1(n593), .B2(\dp/a_neg_mult_id_exe_int[1] ), .A(
        \dp/b10_1_mult_id_exe_int[1] ), .ZN(n5713) );
  OAI211_X1 U6469 ( .C1(\dp/a_mult_id_exe_int[2] ), .C2(n5169), .A(n5711), .B(
        n5710), .ZN(n5816) );
  NAND2_X1 U6470 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[2] ), .A2(n5187), .ZN(
        n5710) );
  NAND2_X1 U6471 ( .A1(\dp/exs/alu_unit/mult/neg_a_shiftn[2] ), .A2(n5188), 
        .ZN(n5711) );
  NOR2_X1 U6472 ( .A1(n5709), .A2(n5708), .ZN(n5719) );
  OAI22_X1 U6473 ( .A1(n5151), .A2(n4105), .B1(n3944), .B2(n4071), .ZN(n5708)
         );
  OAI22_X1 U6474 ( .A1(n3960), .A2(n4227), .B1(n3951), .B2(n4108), .ZN(n5709)
         );
  NOR2_X1 U6475 ( .A1(n3900), .A2(\dp/a_mult_id_exe_int[4] ), .ZN(n5703) );
  NOR2_X1 U6476 ( .A1(n3900), .A2(\dp/a_mult_id_exe_int[3] ), .ZN(n5702) );
  NOR2_X1 U6477 ( .A1(n5696), .A2(n5695), .ZN(n5872) );
  OAI22_X1 U6478 ( .A1(n3960), .A2(n4105), .B1(n3944), .B2(n6459), .ZN(n5695)
         );
  OAI22_X1 U6479 ( .A1(n5151), .A2(n4104), .B1(n3951), .B2(n4223), .ZN(n5696)
         );
  NOR2_X1 U6480 ( .A1(n3900), .A2(\dp/a_mult_id_exe_int[5] ), .ZN(n5692) );
  NOR2_X1 U6481 ( .A1(n3900), .A2(\dp/a_mult_id_exe_int[6] ), .ZN(n5689) );
  OR2_X1 U6482 ( .A1(n5925), .A2(n5089), .ZN(n5090) );
  NOR2_X1 U6483 ( .A1(n5169), .A2(\dp/a_mult_id_exe_int[11] ), .ZN(n5740) );
  OAI211_X1 U6484 ( .C1(n6328), .C2(n6043), .A(n6042), .B(n6041), .ZN(n6056)
         );
  AOI22_X1 U6485 ( .A1(\dp/exs/alu_unit/mult/a_shiftn[24] ), .A2(n3945), .B1(
        n6327), .B2(n4284), .ZN(n6041) );
  AOI22_X1 U6486 ( .A1(n5188), .A2(\dp/exs/alu_unit/mult/neg_a_shiftn[24] ), 
        .B1(\dp/exs/alu_unit/mult/neg_a_shiftn[23] ), .B2(n5154), .ZN(n6042)
         );
  XNOR2_X1 U6487 ( .A(n5146), .B(n5147), .ZN(n5685) );
  INV_X1 U6488 ( .A(\dp/exs/alu_unit/mult/a_shiftn[23] ), .ZN(n6043) );
  OAI211_X1 U6489 ( .C1(n3930), .C2(n4084), .A(n6045), .B(n6044), .ZN(n6057)
         );
  NAND2_X1 U6490 ( .A1(n3943), .A2(\dp/a_neg_mult_id_exe_int[23] ), .ZN(n6044)
         );
  AND2_X1 U6491 ( .A1(n3899), .A2(\dp/b10_1_mult_id_exe_int[1] ), .ZN(n5682)
         );
  AND2_X1 U6492 ( .A1(n6176), .A2(n6178), .ZN(n4873) );
  INV_X1 U6493 ( .A(n7108), .ZN(n6402) );
  NAND2_X1 U6494 ( .A1(n6177), .A2(predicted_taken), .ZN(n4874) );
  NOR2_X1 U6495 ( .A1(n4444), .A2(\ctrl_u/curr_exe[19] ), .ZN(n5823) );
  OAI22_X1 U6496 ( .A1(\dp/npc_id_exe_int[23] ), .A2(\dp/imm_id_exe_int[23] ), 
        .B1(n4275), .B2(n4823), .ZN(n4822) );
  INV_X1 U6497 ( .A(n4827), .ZN(n4823) );
  OAI21_X1 U6498 ( .B1(n4847), .B2(n4828), .A(n4846), .ZN(n4827) );
  NAND2_X1 U6499 ( .A1(n4103), .A2(n4220), .ZN(n4846) );
  NAND2_X1 U6500 ( .A1(n4101), .A2(n4222), .ZN(n4828) );
  NAND2_X1 U6501 ( .A1(n4824), .A2(n4122), .ZN(n4747) );
  NOR2_X1 U6502 ( .A1(n4275), .A2(n4825), .ZN(n4824) );
  INV_X1 U6503 ( .A(n4829), .ZN(n4825) );
  NOR2_X1 U6504 ( .A1(n4830), .A2(n4847), .ZN(n4829) );
  NOR2_X1 U6505 ( .A1(n4103), .A2(n4220), .ZN(n4847) );
  INV_X1 U6506 ( .A(n4941), .ZN(n4830) );
  OAI22_X1 U6507 ( .A1(\dp/npc_id_exe_int[17] ), .A2(n4115), .B1(n4276), .B2(
        n4925), .ZN(n4924) );
  INV_X1 U6508 ( .A(n4929), .ZN(n4925) );
  OAI21_X1 U6509 ( .B1(n4947), .B2(n4930), .A(n4946), .ZN(n4929) );
  NAND2_X1 U6510 ( .A1(n4102), .A2(n4219), .ZN(n4946) );
  NAND2_X1 U6511 ( .A1(n4207), .A2(n4070), .ZN(n4930) );
  NOR2_X1 U6512 ( .A1(n4276), .A2(n4927), .ZN(n4926) );
  INV_X1 U6513 ( .A(n4931), .ZN(n4927) );
  NOR2_X1 U6514 ( .A1(n4932), .A2(n4947), .ZN(n4931) );
  NOR2_X1 U6515 ( .A1(n4102), .A2(n4219), .ZN(n4947) );
  INV_X1 U6516 ( .A(n5002), .ZN(n4932) );
  INV_X1 U6517 ( .A(n5072), .ZN(n5041) );
  INV_X1 U6518 ( .A(n5082), .ZN(n5057) );
  OAI22_X1 U6519 ( .A1(n4048), .A2(n6821), .B1(n4051), .B2(n633), .ZN(n2958)
         );
  OAI22_X1 U6520 ( .A1(n7058), .A2(n6862), .B1(n4049), .B2(n620), .ZN(n2971)
         );
  OAI22_X1 U6521 ( .A1(n4048), .A2(n6782), .B1(n4051), .B2(n640), .ZN(n2951)
         );
  AOI21_X1 U6522 ( .B1(\dp/ids/rp1[27] ), .B2(n4136), .A(n6777), .ZN(n6782) );
  NOR2_X1 U6523 ( .A1(n5230), .A2(n385), .ZN(n6777) );
  OAI22_X1 U6524 ( .A1(n4047), .A2(n6857), .B1(n4050), .B2(n621), .ZN(n2970)
         );
  OAI22_X1 U6525 ( .A1(n4048), .A2(n6826), .B1(n4051), .B2(n632), .ZN(n2959)
         );
  OAI22_X1 U6526 ( .A1(n7058), .A2(n6879), .B1(n4049), .B2(n617), .ZN(n2974)
         );
  AOI21_X1 U6527 ( .B1(\dp/ids/rp1[4] ), .B2(n4136), .A(n6874), .ZN(n6879) );
  NOR2_X1 U6528 ( .A1(n4136), .A2(n362), .ZN(n6874) );
  OAI22_X1 U6529 ( .A1(n7058), .A2(n6882), .B1(n4049), .B2(n616), .ZN(n2975)
         );
  AOI21_X1 U6530 ( .B1(\dp/ids/rp1[3] ), .B2(n4136), .A(n6880), .ZN(n6882) );
  NOR2_X1 U6531 ( .A1(n4136), .A2(n361), .ZN(n6880) );
  OAI22_X1 U6532 ( .A1(n4047), .A2(n6806), .B1(n4050), .B2(n636), .ZN(n2955)
         );
  AOI21_X1 U6533 ( .B1(\dp/ids/rp1[23] ), .B2(n4136), .A(n6801), .ZN(n6806) );
  NOR2_X1 U6534 ( .A1(n5230), .A2(n381), .ZN(n6801) );
  OAI22_X1 U6535 ( .A1(n4047), .A2(n6851), .B1(n4050), .B2(n624), .ZN(n2967)
         );
  OAI22_X1 U6536 ( .A1(n4048), .A2(n6800), .B1(n4051), .B2(n637), .ZN(n2954)
         );
  AOI21_X1 U6537 ( .B1(\dp/ids/rp1[24] ), .B2(n4136), .A(n6795), .ZN(n6800) );
  NOR2_X1 U6538 ( .A1(n5230), .A2(n382), .ZN(n6795) );
  OAI22_X1 U6539 ( .A1(n7058), .A2(n6776), .B1(n4049), .B2(n641), .ZN(n2950)
         );
  AOI21_X1 U6540 ( .B1(\dp/ids/rp1[28] ), .B2(n4136), .A(n6771), .ZN(n6776) );
  NOR2_X1 U6541 ( .A1(n5230), .A2(n386), .ZN(n6771) );
  OAI22_X1 U6542 ( .A1(n4048), .A2(n6849), .B1(n4051), .B2(n625), .ZN(n2966)
         );
  OAI22_X1 U6543 ( .A1(n4050), .A2(n4260), .B1(n4047), .B2(n7042), .ZN(n2717)
         );
  AOI21_X1 U6544 ( .B1(\dp/imm_id_int[4] ), .B2(n4357), .A(n6936), .ZN(n7042)
         );
  NOR2_X1 U6545 ( .A1(n7045), .A2(n4357), .ZN(n6936) );
  OAI22_X1 U6546 ( .A1(n4051), .A2(n4261), .B1(n7058), .B2(n7047), .ZN(n2718)
         );
  AOI21_X1 U6547 ( .B1(\dp/imm_id_int[3] ), .B2(n4357), .A(n6899), .ZN(n7047)
         );
  NOR2_X1 U6548 ( .A1(n7050), .A2(n4357), .ZN(n6899) );
  OAI22_X1 U6549 ( .A1(n4051), .A2(n627), .B1(n4047), .B2(n6844), .ZN(n2964)
         );
  AOI21_X1 U6550 ( .B1(\dp/ids/rp1[14] ), .B2(n4136), .A(n6842), .ZN(n6844) );
  NOR2_X1 U6551 ( .A1(n4136), .A2(n372), .ZN(n6842) );
  OAI22_X1 U6552 ( .A1(n4049), .A2(n631), .B1(n4048), .B2(n6832), .ZN(n2960)
         );
  AOI21_X1 U6553 ( .B1(\dp/ids/rp1[18] ), .B2(n5230), .A(n6827), .ZN(n6832) );
  NOR2_X1 U6554 ( .A1(n5230), .A2(n376), .ZN(n6827) );
  OAI22_X1 U6555 ( .A1(n4050), .A2(n630), .B1(n4048), .B2(n6835), .ZN(n2961)
         );
  AOI21_X1 U6556 ( .B1(\dp/ids/rp1[17] ), .B2(n5230), .A(n6833), .ZN(n6835) );
  NOR2_X1 U6557 ( .A1(n5230), .A2(n375), .ZN(n6833) );
  OAI22_X1 U6558 ( .A1(n4049), .A2(n4264), .B1(n7058), .B2(n7061), .ZN(n2721)
         );
  AOI21_X1 U6559 ( .B1(\dp/ids/rp2[0] ), .B2(b_selector_id), .A(n7055), .ZN(
        n7061) );
  NOR2_X1 U6560 ( .A1(n4477), .A2(b_selector_id), .ZN(n7055) );
  NAND4_X1 U6561 ( .A1(n6958), .A2(n6956), .A3(n6955), .A4(n6954), .ZN(n2695)
         );
  AOI22_X1 U6562 ( .A1(n3898), .A2(\dp/id_exe_regs/b_mult_reg/q[21] ), .B1(
        n3956), .B2(\dp/id_exe_regs/b_mult_reg/q[23] ), .ZN(n6954) );
  OR2_X1 U6563 ( .A1(n4820), .A2(n4603), .ZN(n6955) );
  NAND2_X1 U6564 ( .A1(n5214), .A2(\dp/ids/rp2[22] ), .ZN(n6956) );
  NAND4_X1 U6565 ( .A1(n6958), .A2(n6953), .A3(n6952), .A4(n6951), .ZN(n2699)
         );
  AOI22_X1 U6566 ( .A1(n3897), .A2(\dp/id_exe_regs/b_mult_reg/q[17] ), .B1(
        n3947), .B2(\dp/id_exe_regs/b_mult_reg/q[19] ), .ZN(n6951) );
  NAND2_X1 U6567 ( .A1(n4648), .A2(rt_id[2]), .ZN(n6952) );
  NAND2_X1 U6568 ( .A1(n5214), .A2(\dp/ids/rp2[18] ), .ZN(n6953) );
  AOI22_X1 U6569 ( .A1(n3897), .A2(\dp/id_exe_regs/b_mult_reg/q[23] ), .B1(
        n3956), .B2(\dp/id_exe_regs/b_mult_reg/q[25] ), .ZN(n6957) );
  NAND4_X1 U6570 ( .A1(n6958), .A2(n6918), .A3(n6917), .A4(n6916), .ZN(n2696)
         );
  AOI22_X1 U6571 ( .A1(n3896), .A2(\dp/id_exe_regs/b_mult_reg/q[20] ), .B1(
        n3956), .B2(\dp/id_exe_regs/b_mult_reg/q[22] ), .ZN(n6916) );
  NAND2_X1 U6572 ( .A1(n4648), .A2(rs_id[0]), .ZN(n6917) );
  INV_X1 U6573 ( .A(n7436), .ZN(n6981) );
  NAND2_X1 U6574 ( .A1(n5214), .A2(\dp/ids/rp2[21] ), .ZN(n6918) );
  INV_X1 U6575 ( .A(n4820), .ZN(n6923) );
  NAND2_X1 U6576 ( .A1(n3901), .A2(n4111), .ZN(n4820) );
  OAI211_X1 U6577 ( .C1(n5215), .C2(n6999), .A(n6998), .B(n6997), .ZN(n2739)
         );
  NAND2_X1 U6578 ( .A1(n5216), .A2(n4410), .ZN(n6997) );
  NAND2_X1 U6579 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[17] ), .ZN(n6998) );
  INV_X1 U6580 ( .A(\dp/ids/rp2[17] ), .ZN(n6999) );
  OAI211_X1 U6581 ( .C1(n5215), .C2(n7004), .A(n7003), .B(n7002), .ZN(n2740)
         );
  NAND2_X1 U6582 ( .A1(n5216), .A2(n4411), .ZN(n7002) );
  NAND2_X1 U6583 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[16] ), .ZN(n7003) );
  INV_X1 U6584 ( .A(\dp/ids/rp2[16] ), .ZN(n7004) );
  OAI22_X1 U6585 ( .A1(n4051), .A2(n639), .B1(n7058), .B2(n6788), .ZN(n2952)
         );
  AOI21_X1 U6586 ( .B1(\dp/ids/rp1[26] ), .B2(n4136), .A(n6783), .ZN(n6788) );
  NOR2_X1 U6587 ( .A1(n5230), .A2(n384), .ZN(n6783) );
  OAI22_X1 U6588 ( .A1(n4049), .A2(n622), .B1(n4047), .B2(n6855), .ZN(n2969)
         );
  OAI22_X1 U6589 ( .A1(n4050), .A2(n634), .B1(n4048), .B2(n6816), .ZN(n2957)
         );
  OAI22_X1 U6590 ( .A1(n4050), .A2(n626), .B1(n4047), .B2(n6847), .ZN(n2965)
         );
  AOI21_X1 U6591 ( .B1(\dp/ids/rp1[13] ), .B2(n4136), .A(n6845), .ZN(n6847) );
  NOR2_X1 U6592 ( .A1(n4136), .A2(n371), .ZN(n6845) );
  OAI22_X1 U6593 ( .A1(n4051), .A2(n623), .B1(n7058), .B2(n6853), .ZN(n2968)
         );
  OAI22_X1 U6594 ( .A1(n4051), .A2(n618), .B1(n4047), .B2(n6873), .ZN(n2973)
         );
  OAI22_X1 U6595 ( .A1(n4049), .A2(n619), .B1(n4048), .B2(n6868), .ZN(n2972)
         );
  AOI21_X1 U6596 ( .B1(\dp/ids/rp1[6] ), .B2(n4136), .A(n6863), .ZN(n6868) );
  NOR2_X1 U6597 ( .A1(n4136), .A2(n364), .ZN(n6863) );
  OAI22_X1 U6598 ( .A1(n4050), .A2(n642), .B1(n4048), .B2(n6770), .ZN(n2949)
         );
  AOI21_X1 U6599 ( .B1(\dp/ids/rp1[29] ), .B2(n4136), .A(n6765), .ZN(n6770) );
  NOR2_X1 U6600 ( .A1(n4136), .A2(n387), .ZN(n6765) );
  OAI22_X1 U6601 ( .A1(n4049), .A2(n615), .B1(n7058), .B2(n6884), .ZN(n2976)
         );
  OAI22_X1 U6602 ( .A1(n4051), .A2(n635), .B1(n7058), .B2(n6811), .ZN(n2956)
         );
  OAI22_X1 U6603 ( .A1(n4049), .A2(n643), .B1(n4047), .B2(n6764), .ZN(n2948)
         );
  AOI21_X1 U6604 ( .B1(\dp/ids/rp1[30] ), .B2(n4136), .A(n6759), .ZN(n6764) );
  NOR2_X1 U6605 ( .A1(n5230), .A2(n388), .ZN(n6759) );
  OAI22_X1 U6606 ( .A1(n4050), .A2(n638), .B1(n4048), .B2(n6794), .ZN(n2953)
         );
  AOI21_X1 U6607 ( .B1(\dp/ids/rp1[25] ), .B2(n4136), .A(n6789), .ZN(n6794) );
  NOR2_X1 U6608 ( .A1(n5230), .A2(n383), .ZN(n6789) );
  OAI21_X1 U6609 ( .B1(n3934), .B2(n4544), .A(n5546), .ZN(\ctrl_u/n537 ) );
  AOI211_X1 U6610 ( .C1(n5627), .C2(n5543), .A(n5590), .B(n3962), .ZN(n5544)
         );
  NOR2_X1 U6611 ( .A1(instr_if[28]), .A2(n7275), .ZN(n5552) );
  INV_X1 U6612 ( .A(n5645), .ZN(n5543) );
  NOR2_X1 U6613 ( .A1(instr_if[31]), .A2(n5560), .ZN(n5645) );
  NOR3_X1 U6614 ( .A1(instr_if[2]), .A2(n5542), .A3(n7279), .ZN(n5545) );
  AOI22_X1 U6615 ( .A1(instr_if[1]), .A2(n5541), .B1(instr_if[0]), .B2(n5540), 
        .ZN(n5542) );
  NAND2_X1 U6616 ( .A1(n7029), .A2(n4697), .ZN(n2748) );
  NAND2_X1 U6617 ( .A1(n4682), .A2(\dp/ids/rp2[8] ), .ZN(n4697) );
  AOI22_X1 U6618 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[8] ), .B1(n4107), .B2(
        n4432), .ZN(n7029) );
  NAND2_X1 U6619 ( .A1(n7014), .A2(n4676), .ZN(n2743) );
  NAND2_X1 U6620 ( .A1(n3955), .A2(\dp/ids/rp2[13] ), .ZN(n4676) );
  AOI22_X1 U6621 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[13] ), .B1(n5217), .B2(
        n4427), .ZN(n7014) );
  NAND2_X1 U6622 ( .A1(n7023), .A2(n4677), .ZN(n2746) );
  NAND2_X1 U6623 ( .A1(n3955), .A2(\dp/ids/rp2[10] ), .ZN(n4677) );
  AOI22_X1 U6624 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[10] ), .B1(n4107), .B2(
        n4430), .ZN(n7023) );
  NAND2_X1 U6625 ( .A1(n7020), .A2(n4696), .ZN(n2745) );
  NAND2_X1 U6626 ( .A1(n3955), .A2(\dp/ids/rp2[11] ), .ZN(n4696) );
  AOI22_X1 U6627 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[11] ), .B1(n5217), .B2(
        n4429), .ZN(n7020) );
  NAND2_X1 U6628 ( .A1(n7008), .A2(n4679), .ZN(n2741) );
  NAND2_X1 U6629 ( .A1(n4682), .A2(\dp/ids/rp2[15] ), .ZN(n4679) );
  AOI22_X1 U6630 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[15] ), .B1(n5216), .B2(
        n4425), .ZN(n7008) );
  NAND2_X1 U6631 ( .A1(n7026), .A2(n4681), .ZN(n2747) );
  NAND2_X1 U6632 ( .A1(n4682), .A2(\dp/ids/rp2[9] ), .ZN(n4681) );
  AOI22_X1 U6633 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[9] ), .B1(n5216), .B2(
        n4431), .ZN(n7026) );
  NAND2_X1 U6634 ( .A1(n7035), .A2(n4683), .ZN(n2750) );
  NAND2_X1 U6635 ( .A1(n4682), .A2(\dp/ids/rp2[6] ), .ZN(n4683) );
  AOI22_X1 U6636 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[6] ), .B1(n5217), .B2(
        n4434), .ZN(n7035) );
  NAND2_X1 U6637 ( .A1(n7032), .A2(n4678), .ZN(n2749) );
  NAND2_X1 U6638 ( .A1(n3955), .A2(\dp/ids/rp2[7] ), .ZN(n4678) );
  AOI22_X1 U6639 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[7] ), .B1(n5216), .B2(
        n4433), .ZN(n7032) );
  NAND2_X1 U6640 ( .A1(n7040), .A2(n4698), .ZN(n2751) );
  NAND2_X1 U6641 ( .A1(n3955), .A2(\dp/ids/rp2[5] ), .ZN(n4698) );
  AOI22_X1 U6642 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[5] ), .B1(n5217), .B2(
        n4435), .ZN(n7040) );
  NAND2_X1 U6643 ( .A1(n7017), .A2(n4680), .ZN(n2744) );
  NAND2_X1 U6644 ( .A1(n4682), .A2(\dp/ids/rp2[12] ), .ZN(n4680) );
  AND2_X1 U6645 ( .A1(n3902), .A2(n4584), .ZN(n6930) );
  AOI22_X1 U6646 ( .A1(n5129), .A2(\dp/op_b_id_ex_int[12] ), .B1(n5217), .B2(
        n4428), .ZN(n7017) );
  AND4_X1 U6647 ( .A1(n5500), .A2(n5499), .A3(n5596), .A4(n7277), .ZN(n5534)
         );
  NOR2_X1 U6648 ( .A1(instr_if[4]), .A2(n5497), .ZN(n5500) );
  NAND2_X1 U6649 ( .A1(n3948), .A2(n5339), .ZN(n4965) );
  OAI22_X1 U6650 ( .A1(instr_if[26]), .A2(n5532), .B1(n5531), .B2(n5530), .ZN(
        n5533) );
  NAND2_X1 U6651 ( .A1(n7264), .A2(n5540), .ZN(n5531) );
  INV_X1 U6652 ( .A(n5519), .ZN(n5540) );
  INV_X1 U6653 ( .A(n5529), .ZN(n5532) );
  NOR2_X1 U6654 ( .A1(instr_if[31]), .A2(n5522), .ZN(n5529) );
  INV_X1 U6655 ( .A(n5528), .ZN(n5536) );
  AOI21_X1 U6656 ( .B1(n5591), .B2(n5520), .A(n5524), .ZN(n5521) );
  NOR3_X1 U6657 ( .A1(n5530), .A2(n5519), .A3(n5518), .ZN(n5524) );
  NAND2_X1 U6658 ( .A1(n7280), .A2(n7279), .ZN(n5518) );
  NAND2_X1 U6659 ( .A1(n5541), .A2(n7278), .ZN(n5519) );
  NOR3_X1 U6660 ( .A1(n5594), .A2(n5497), .A3(n7277), .ZN(n5541) );
  INV_X1 U6661 ( .A(n7293), .ZN(n5497) );
  INV_X1 U6662 ( .A(n5499), .ZN(n5594) );
  INV_X1 U6663 ( .A(n5522), .ZN(n5520) );
  INV_X1 U6664 ( .A(n5506), .ZN(n5591) );
  NAND2_X1 U6665 ( .A1(n5627), .A2(n5644), .ZN(n5506) );
  OR2_X1 U6666 ( .A1(n4968), .A2(\ctrl_u/if_stall ), .ZN(n4854) );
  INV_X1 U6667 ( .A(n5176), .ZN(n4651) );
  OAI22_X1 U6668 ( .A1(n5458), .A2(n5457), .B1(\ctrl_u/curr_id[34] ), .B2(
        n5599), .ZN(n4667) );
  OAI21_X1 U6669 ( .B1(n5491), .B2(n5514), .A(n5456), .ZN(n5457) );
  NAND2_X1 U6670 ( .A1(instr_if[29]), .A2(instr_if[30]), .ZN(n5491) );
  OAI22_X1 U6671 ( .A1(n5458), .A2(n5436), .B1(\ctrl_u/curr_id[35] ), .B2(
        n5599), .ZN(n4674) );
  OAI22_X1 U6672 ( .A1(n7291), .A2(n5483), .B1(n5589), .B2(n5630), .ZN(n5436)
         );
  NAND2_X1 U6673 ( .A1(instr_if[28]), .A2(instr_if[30]), .ZN(n5630) );
  INV_X1 U6674 ( .A(n5490), .ZN(n5589) );
  NAND2_X1 U6675 ( .A1(n5499), .A2(n7264), .ZN(n5483) );
  NAND2_X1 U6676 ( .A1(n5016), .A2(n5015), .ZN(n5458) );
  AND3_X1 U6677 ( .A1(n5435), .A2(n5465), .A3(n5434), .ZN(n5015) );
  NAND2_X1 U6678 ( .A1(n5499), .A2(n5433), .ZN(n5434) );
  OAI211_X1 U6679 ( .C1(n7264), .C2(n7285), .A(n7286), .B(n5432), .ZN(n5433)
         );
  AOI22_X1 U6680 ( .A1(n7287), .A2(n7288), .B1(n5501), .B2(n5455), .ZN(n5432)
         );
  INV_X1 U6681 ( .A(n7291), .ZN(n5455) );
  NOR2_X1 U6682 ( .A1(n7279), .A2(n7281), .ZN(n5501) );
  INV_X1 U6683 ( .A(instr_if[4]), .ZN(n7278) );
  NAND2_X1 U6684 ( .A1(n7280), .A2(n5530), .ZN(n7284) );
  NAND2_X1 U6685 ( .A1(instr_if[5]), .A2(n5596), .ZN(n7285) );
  NOR2_X1 U6686 ( .A1(n7280), .A2(n5530), .ZN(n5596) );
  NOR2_X1 U6687 ( .A1(instr_if[3]), .A2(instr_if[0]), .ZN(n7264) );
  NOR2_X1 U6688 ( .A1(instr_if[26]), .A2(n5502), .ZN(n5499) );
  NAND2_X1 U6689 ( .A1(n5427), .A2(n5627), .ZN(n5502) );
  NAND2_X1 U6690 ( .A1(instr_if[31]), .A2(n5648), .ZN(n5465) );
  NAND2_X1 U6691 ( .A1(n5647), .A2(n5504), .ZN(n5435) );
  NOR2_X1 U6692 ( .A1(n5648), .A2(n5494), .ZN(n5504) );
  NOR2_X1 U6693 ( .A1(instr_if[29]), .A2(n5590), .ZN(n5647) );
  NOR2_X1 U6694 ( .A1(n5626), .A2(n5017), .ZN(n5016) );
  OR3_X1 U6695 ( .A1(n5643), .A2(n5431), .A3(n5637), .ZN(n5017) );
  NOR2_X1 U6696 ( .A1(n5496), .A2(n5450), .ZN(n5637) );
  INV_X1 U6697 ( .A(n5638), .ZN(n5450) );
  NOR2_X1 U6698 ( .A1(n5430), .A2(n5562), .ZN(n5638) );
  NAND2_X1 U6699 ( .A1(instr_if[26]), .A2(n5627), .ZN(n5562) );
  INV_X1 U6700 ( .A(n5427), .ZN(n5430) );
  NOR2_X1 U6701 ( .A1(instr_if[28]), .A2(n5651), .ZN(n5427) );
  NAND2_X1 U6702 ( .A1(n5445), .A2(n5590), .ZN(n5651) );
  NOR2_X1 U6703 ( .A1(instr_if[29]), .A2(instr_if[31]), .ZN(n5445) );
  NOR4_X1 U6704 ( .A1(instr_if[20]), .A2(instr_if[19]), .A3(instr_if[18]), 
        .A4(instr_if[17]), .ZN(n5496) );
  NOR3_X1 U6705 ( .A1(n5560), .A2(n5514), .A3(n7275), .ZN(n5431) );
  INV_X1 U6706 ( .A(n5648), .ZN(n5514) );
  NOR2_X1 U6707 ( .A1(n5627), .A2(n7276), .ZN(n5648) );
  INV_X1 U6708 ( .A(instr_if[28]), .ZN(n7276) );
  OAI21_X1 U6709 ( .B1(n5644), .B2(n5522), .A(n5475), .ZN(n5643) );
  AOI22_X1 U6710 ( .A1(n5553), .A2(n5490), .B1(instr_if[30]), .B2(n5440), .ZN(
        n5475) );
  INV_X1 U6711 ( .A(n5633), .ZN(n5440) );
  NAND2_X1 U6712 ( .A1(instr_if[31]), .A2(n5494), .ZN(n5633) );
  NOR2_X1 U6713 ( .A1(instr_if[27]), .A2(instr_if[28]), .ZN(n5494) );
  NOR2_X1 U6714 ( .A1(instr_if[26]), .A2(n5627), .ZN(n5490) );
  INV_X1 U6715 ( .A(n5548), .ZN(n5553) );
  NAND2_X1 U6716 ( .A1(instr_if[31]), .A2(n5590), .ZN(n5548) );
  NAND2_X1 U6717 ( .A1(n5419), .A2(n4237), .ZN(n5421) );
  NAND2_X1 U6718 ( .A1(n5659), .A2(n5618), .ZN(n5419) );
  NAND2_X1 U6719 ( .A1(n5675), .A2(n5097), .ZN(n5659) );
  NAND2_X1 U6720 ( .A1(n5422), .A2(\ctrl_u/n555 ), .ZN(n4966) );
  NOR2_X1 U6721 ( .A1(n4237), .A2(n7340), .ZN(n5418) );
  AOI21_X1 U6722 ( .B1(n5341), .B2(n5340), .A(n4303), .ZN(n5675) );
  NAND4_X1 U6723 ( .A1(n4736), .A2(n4737), .A3(n3909), .A4(n4959), .ZN(n5341)
         );
  NAND2_X1 U6724 ( .A1(n4056), .A2(n6749), .ZN(n2889) );
  NAND2_X1 U6725 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[57] ), .ZN(n6749) );
  NAND2_X1 U6726 ( .A1(n4055), .A2(n6740), .ZN(n2898) );
  NAND2_X1 U6727 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[48] ), .ZN(n6740) );
  NAND2_X1 U6728 ( .A1(n4056), .A2(n6733), .ZN(n2905) );
  NAND2_X1 U6729 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[41] ), .ZN(n6733) );
  NAND2_X1 U6730 ( .A1(n4057), .A2(n6747), .ZN(n2891) );
  NAND2_X1 U6731 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[55] ), .ZN(n6747) );
  NAND2_X1 U6732 ( .A1(n4056), .A2(n6746), .ZN(n2892) );
  NAND2_X1 U6733 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[54] ), .ZN(n6746) );
  NAND2_X1 U6734 ( .A1(n4055), .A2(n6745), .ZN(n2893) );
  NAND2_X1 U6735 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[53] ), .ZN(n6745) );
  NAND2_X1 U6736 ( .A1(n4055), .A2(n6731), .ZN(n2907) );
  NAND2_X1 U6737 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[39] ), .ZN(n6731) );
  NAND2_X1 U6738 ( .A1(n4056), .A2(n6728), .ZN(n2910) );
  NAND2_X1 U6739 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[36] ), .ZN(n6728) );
  NAND2_X1 U6740 ( .A1(n4057), .A2(n6755), .ZN(n2883) );
  NAND2_X1 U6741 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[63] ), .ZN(n6755) );
  NAND2_X1 U6742 ( .A1(n4056), .A2(n6738), .ZN(n2900) );
  NAND2_X1 U6743 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[46] ), .ZN(n6738) );
  NAND2_X1 U6744 ( .A1(n4056), .A2(n6743), .ZN(n2895) );
  NAND2_X1 U6745 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[51] ), .ZN(n6743) );
  NAND2_X1 U6746 ( .A1(n4056), .A2(n6742), .ZN(n2896) );
  NAND2_X1 U6747 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[50] ), .ZN(n6742) );
  NAND2_X1 U6748 ( .A1(n4057), .A2(n6734), .ZN(n2904) );
  NAND2_X1 U6749 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[42] ), .ZN(n6734) );
  NAND2_X1 U6750 ( .A1(n4055), .A2(n6744), .ZN(n2894) );
  NAND2_X1 U6751 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[52] ), .ZN(n6744) );
  NAND2_X1 U6752 ( .A1(n4057), .A2(n6741), .ZN(n2897) );
  NAND2_X1 U6753 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[49] ), .ZN(n6741) );
  NAND2_X1 U6754 ( .A1(n4057), .A2(n6735), .ZN(n2903) );
  NAND2_X1 U6755 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[43] ), .ZN(n6735) );
  NAND2_X1 U6756 ( .A1(n4056), .A2(n6739), .ZN(n2899) );
  NAND2_X1 U6757 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[47] ), .ZN(n6739) );
  NAND2_X1 U6758 ( .A1(n4055), .A2(n6732), .ZN(n2906) );
  NAND2_X1 U6759 ( .A1(n3877), .A2(\dp/a_mult_id_exe_int[40] ), .ZN(n6732) );
  NAND2_X1 U6760 ( .A1(n4056), .A2(n6729), .ZN(n2909) );
  NAND2_X1 U6761 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[37] ), .ZN(n6729) );
  NAND2_X1 U6762 ( .A1(n4056), .A2(n6737), .ZN(n2901) );
  NAND2_X1 U6763 ( .A1(n3876), .A2(\dp/a_mult_id_exe_int[45] ), .ZN(n6737) );
  NAND2_X1 U6764 ( .A1(n4055), .A2(n6730), .ZN(n2908) );
  NAND2_X1 U6765 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[38] ), .ZN(n6730) );
  NAND2_X1 U6766 ( .A1(n4057), .A2(n6736), .ZN(n2902) );
  NAND2_X1 U6767 ( .A1(n3878), .A2(\dp/a_mult_id_exe_int[44] ), .ZN(n6736) );
  NAND2_X1 U6768 ( .A1(n6472), .A2(n6471), .ZN(n6722) );
  NAND2_X1 U6769 ( .A1(n4358), .A2(n4384), .ZN(n6471) );
  NAND2_X1 U6770 ( .A1(\dp/ids/rp1[31] ), .A2(n4136), .ZN(n6472) );
  INV_X1 U6771 ( .A(n6721), .ZN(n4914) );
  NAND4_X1 U6772 ( .A1(n7310), .A2(n7311), .A3(n5388), .A4(n5387), .ZN(n7312)
         );
  NAND2_X1 U6773 ( .A1(n5386), .A2(\ctrl_u/curr_wb[3] ), .ZN(n5387) );
  OAI22_X1 U6774 ( .A1(n5385), .A2(n5384), .B1(n5383), .B2(n5382), .ZN(n5386)
         );
  NAND2_X1 U6775 ( .A1(n5381), .A2(n5380), .ZN(n5382) );
  XNOR2_X1 U6776 ( .A(rs_id[1]), .B(rd[1]), .ZN(n5380) );
  XNOR2_X1 U6777 ( .A(rs_id[3]), .B(rd[3]), .ZN(n5381) );
  XNOR2_X1 U6778 ( .A(rs_id[2]), .B(rd[2]), .ZN(n5377) );
  XNOR2_X1 U6779 ( .A(rs_id[4]), .B(rd[4]), .ZN(n5378) );
  AOI21_X1 U6780 ( .B1(n4083), .B2(rd[0]), .A(n5376), .ZN(n5379) );
  NOR2_X1 U6781 ( .A1(rd[0]), .A2(n4083), .ZN(n5376) );
  XNOR2_X1 U6782 ( .A(rt_id[2]), .B(rd[2]), .ZN(n5373) );
  XNOR2_X1 U6783 ( .A(rt_id[0]), .B(rd[0]), .ZN(n5374) );
  AOI21_X1 U6784 ( .B1(n4212), .B2(rd[3]), .A(n5372), .ZN(n5375) );
  NOR2_X1 U6785 ( .A1(rd[3]), .A2(n4212), .ZN(n5372) );
  NAND2_X1 U6786 ( .A1(n5371), .A2(n5370), .ZN(n5385) );
  XNOR2_X1 U6787 ( .A(rt_id[1]), .B(rd[1]), .ZN(n5370) );
  XNOR2_X1 U6788 ( .A(rt_id[4]), .B(rd[4]), .ZN(n5371) );
  AOI21_X1 U6789 ( .B1(n4299), .B2(n7309), .A(n5369), .ZN(n5388) );
  NOR2_X1 U6790 ( .A1(n5368), .A2(n5367), .ZN(n5369) );
  NAND2_X1 U6791 ( .A1(n5366), .A2(n5365), .ZN(n5367) );
  XNOR2_X1 U6792 ( .A(rt_id[1]), .B(n3970), .ZN(n5365) );
  NAND4_X1 U6793 ( .A1(n5364), .A2(\ctrl_u/curr_mem[3] ), .A3(n5363), .A4(
        n5362), .ZN(n5368) );
  XNOR2_X1 U6794 ( .A(rd_exemem[2]), .B(rt_id[2]), .ZN(n5362) );
  XNOR2_X1 U6795 ( .A(n4021), .B(rt_id[4]), .ZN(n5363) );
  XNOR2_X1 U6796 ( .A(rt_id[3]), .B(rd_exemem[3]), .ZN(n5364) );
  XNOR2_X1 U6797 ( .A(n4010), .B(rs_id[3]), .ZN(n5358) );
  XNOR2_X1 U6798 ( .A(rs_id[1]), .B(n3970), .ZN(n5359) );
  XNOR2_X1 U6799 ( .A(rs_id[4]), .B(n4021), .ZN(n5360) );
  NOR2_X1 U6800 ( .A1(n5357), .A2(n4265), .ZN(n5361) );
  NOR2_X1 U6801 ( .A1(n5332), .A2(n4287), .ZN(n5049) );
  NAND2_X1 U6802 ( .A1(n5334), .A2(n6161), .ZN(n6163) );
  INV_X1 U6803 ( .A(n6162), .ZN(n5334) );
  INV_X1 U6804 ( .A(n6161), .ZN(n6159) );
  INV_X1 U6805 ( .A(n4753), .ZN(n4752) );
  NAND2_X1 U6806 ( .A1(n4755), .A2(n4751), .ZN(n4754) );
  INV_X1 U6807 ( .A(n4759), .ZN(n4755) );
  XNOR2_X1 U6808 ( .A(\intadd_1/A[26] ), .B(\intadd_1/B[26] ), .ZN(n4777) );
  INV_X1 U6809 ( .A(n4709), .ZN(n5076) );
  XNOR2_X1 U6810 ( .A(n4729), .B(\intadd_1/n17 ), .ZN(\intadd_1/SUM[9] ) );
  NOR2_X1 U6811 ( .A1(n5001), .A2(n4796), .ZN(n4788) );
  INV_X1 U6812 ( .A(n5001), .ZN(n4789) );
  XNOR2_X1 U6813 ( .A(\intadd_1/A[28] ), .B(\intadd_1/B[28] ), .ZN(n5001) );
  XNOR2_X1 U6814 ( .A(\intadd_1/n104 ), .B(\intadd_1/n13 ), .ZN(
        \intadd_1/SUM[13] ) );
  INV_X1 U6815 ( .A(n4750), .ZN(n4756) );
  OAI21_X1 U6816 ( .B1(n5060), .B2(n4758), .A(n4757), .ZN(n4750) );
  XNOR2_X1 U6817 ( .A(\intadd_1/A[27] ), .B(\intadd_1/B[27] ), .ZN(n4804) );
  XNOR2_X1 U6818 ( .A(\intadd_1/n147 ), .B(\intadd_1/n20 ), .ZN(
        \intadd_1/SUM[6] ) );
  AND3_X1 U6819 ( .A1(\intadd_1/SUM[1] ), .A2(n7067), .A3(\intadd_1/SUM[0] ), 
        .ZN(n5329) );
  AND2_X1 U6820 ( .A1(n7079), .A2(n5328), .ZN(n7067) );
  XNOR2_X1 U6821 ( .A(\intadd_1/n117 ), .B(\intadd_1/n15 ), .ZN(
        \intadd_1/SUM[11] ) );
  OAI21_X1 U6822 ( .B1(\intadd_1/n139 ), .B2(\intadd_1/n118 ), .A(n4027), .ZN(
        \intadd_1/n117 ) );
  INV_X1 U6823 ( .A(n4986), .ZN(n4961) );
  NOR2_X1 U6824 ( .A1(n5048), .A2(n5070), .ZN(n4987) );
  INV_X1 U6825 ( .A(n5332), .ZN(n5048) );
  INV_X1 U6826 ( .A(n5049), .ZN(n4988) );
  XNOR2_X1 U6827 ( .A(n6161), .B(n4225), .ZN(n5333) );
  XNOR2_X1 U6828 ( .A(\intadd_1/n28 ), .B(n5071), .ZN(\intadd_1/SUM[29] ) );
  XNOR2_X1 U6829 ( .A(\intadd_1/A[29] ), .B(\intadd_1/B[29] ), .ZN(n5071) );
  NAND2_X1 U6830 ( .A1(n5280), .A2(n5279), .ZN(n7193) );
  NOR2_X1 U6831 ( .A1(n5175), .A2(n492), .ZN(n5281) );
  INV_X1 U6832 ( .A(wp_data[29]), .ZN(n5278) );
  NOR2_X1 U6833 ( .A1(n5175), .A2(n491), .ZN(n5283) );
  INV_X1 U6834 ( .A(wp_data[28]), .ZN(n5282) );
  NAND2_X1 U6835 ( .A1(\intadd_1/B[22] ), .A2(n4699), .ZN(\intadd_1/n54 ) );
  NAND2_X1 U6836 ( .A1(n4845), .A2(\intadd_1/B[20] ), .ZN(\intadd_1/n62 ) );
  NAND2_X1 U6837 ( .A1(\intadd_1/A[16] ), .A2(\intadd_1/B[16] ), .ZN(
        \intadd_1/n83 ) );
  AOI21_X1 U6838 ( .B1(n5118), .B2(n4243), .A(n7203), .ZN(\intadd_1/B[23] ) );
  INV_X1 U6839 ( .A(wp_data[24]), .ZN(n5288) );
  OAI22_X1 U6840 ( .A1(n5293), .A2(n3950), .B1(n5173), .B2(n4075), .ZN(n7213)
         );
  INV_X1 U6841 ( .A(wp_data[19]), .ZN(n5293) );
  INV_X1 U6842 ( .A(wp_data[18]), .ZN(n5294) );
  NAND2_X1 U6843 ( .A1(n5297), .A2(n5296), .ZN(n7217) );
  OR2_X1 U6844 ( .A1(n5173), .A2(n4095), .ZN(n5297) );
  NOR2_X1 U6845 ( .A1(n3949), .A2(n480), .ZN(n5298) );
  INV_X1 U6846 ( .A(wp_data[17]), .ZN(n5295) );
  NOR2_X1 U6847 ( .A1(n3949), .A2(n479), .ZN(n5300) );
  INV_X1 U6848 ( .A(wp_data[16]), .ZN(n5299) );
  AOI21_X1 U6849 ( .B1(n5118), .B2(n4244), .A(n7205), .ZN(\intadd_1/B[22] ) );
  OAI22_X1 U6850 ( .A1(n5289), .A2(n5172), .B1(n5173), .B2(n4078), .ZN(n7205)
         );
  INV_X1 U6851 ( .A(wp_data[23]), .ZN(n5289) );
  OAI22_X1 U6852 ( .A1(n5290), .A2(n3950), .B1(n5173), .B2(n4077), .ZN(n7207)
         );
  INV_X1 U6853 ( .A(wp_data[22]), .ZN(n5290) );
  AOI21_X1 U6854 ( .B1(n5118), .B2(n4246), .A(n7209), .ZN(\intadd_1/B[20] ) );
  INV_X1 U6855 ( .A(wp_data[21]), .ZN(n5291) );
  OAI22_X1 U6856 ( .A1(n5292), .A2(n5172), .B1(n5173), .B2(n4076), .ZN(n7211)
         );
  INV_X1 U6857 ( .A(wp_data[20]), .ZN(n5292) );
  NAND2_X1 U6858 ( .A1(\intadd_1/A[6] ), .A2(\intadd_1/B[6] ), .ZN(
        \intadd_1/n146 ) );
  NAND2_X1 U6859 ( .A1(n4668), .A2(\intadd_1/B[4] ), .ZN(\intadd_1/n154 ) );
  OAI21_X1 U6860 ( .B1(n5123), .B2(n4377), .A(n5053), .ZN(n7251) );
  NAND2_X1 U6861 ( .A1(n5330), .A2(wp_data[0]), .ZN(n5053) );
  NAND2_X1 U6862 ( .A1(n7259), .A2(n5326), .ZN(n7071) );
  AOI21_X1 U6863 ( .B1(n5325), .B2(n4255), .A(n7249), .ZN(\intadd_1/B[0] ) );
  OAI22_X1 U6864 ( .A1(n5324), .A2(n3950), .B1(n5173), .B2(n4072), .ZN(n7249)
         );
  AND2_X1 U6865 ( .A1(n5119), .A2(\dp/b_adder_id_exe_int[1] ), .ZN(n4733) );
  INV_X1 U6866 ( .A(wp_data[1]), .ZN(n5324) );
  NOR2_X1 U6867 ( .A1(n5175), .A2(n465), .ZN(n5272) );
  OAI22_X1 U6868 ( .A1(n5123), .A2(n4080), .B1(n5321), .B2(n3950), .ZN(n7245)
         );
  INV_X1 U6869 ( .A(wp_data[3]), .ZN(n5321) );
  NOR2_X1 U6870 ( .A1(n3949), .A2(n466), .ZN(n5322) );
  INV_X1 U6871 ( .A(wp_data[6]), .ZN(n5317) );
  OAI22_X1 U6872 ( .A1(n5316), .A2(n3950), .B1(n5173), .B2(n6453), .ZN(n7237)
         );
  INV_X1 U6873 ( .A(wp_data[7]), .ZN(n5316) );
  INV_X1 U6874 ( .A(wp_data[4]), .ZN(n5319) );
  NOR2_X1 U6875 ( .A1(n5174), .A2(n467), .ZN(n5320) );
  NAND2_X1 U6876 ( .A1(n4024), .A2(wp_data[4]), .ZN(n5261) );
  OAI22_X1 U6877 ( .A1(n5318), .A2(n5172), .B1(n5173), .B2(n6459), .ZN(n7241)
         );
  INV_X1 U6878 ( .A(wp_data[5]), .ZN(n5318) );
  NOR2_X1 U6879 ( .A1(n3949), .A2(n478), .ZN(n5302) );
  INV_X1 U6880 ( .A(wp_data[15]), .ZN(n5301) );
  OAI22_X1 U6881 ( .A1(n5303), .A2(n5172), .B1(n5173), .B2(n4066), .ZN(n7223)
         );
  INV_X1 U6882 ( .A(wp_data[14]), .ZN(n5303) );
  OAI22_X1 U6883 ( .A1(n5173), .A2(n4079), .B1(n5304), .B2(n5171), .ZN(n7225)
         );
  INV_X1 U6884 ( .A(wp_data[13]), .ZN(n5304) );
  INV_X1 U6885 ( .A(wp_data[12]), .ZN(n5305) );
  NOR2_X1 U6886 ( .A1(n3949), .A2(n472), .ZN(n5313) );
  NOR2_X1 U6887 ( .A1(n5174), .A2(n471), .ZN(n5315) );
  INV_X1 U6888 ( .A(wp_data[8]), .ZN(n5314) );
  NOR2_X1 U6889 ( .A1(n5175), .A2(n474), .ZN(n5309) );
  OR2_X1 U6890 ( .A1(n5173), .A2(n4073), .ZN(n5308) );
  INV_X1 U6891 ( .A(wp_data[11]), .ZN(n5306) );
  NOR2_X1 U6892 ( .A1(n3949), .A2(n473), .ZN(n5311) );
  INV_X1 U6893 ( .A(wp_data[10]), .ZN(n5310) );
  OAI22_X1 U6894 ( .A1(n4065), .A2(n5173), .B1(n5172), .B2(n5286), .ZN(n7199)
         );
  INV_X1 U6895 ( .A(wp_data[26]), .ZN(n5286) );
  NOR2_X1 U6896 ( .A1(n5174), .A2(n490), .ZN(n5285) );
  INV_X1 U6897 ( .A(wp_data[27]), .ZN(n5284) );
  OAI22_X1 U6898 ( .A1(n4062), .A2(n5173), .B1(n3950), .B2(n5287), .ZN(n7201)
         );
  INV_X1 U6899 ( .A(wp_data[25]), .ZN(n5287) );
  NAND2_X1 U6900 ( .A1(n5086), .A2(n5081), .ZN(n4798) );
  XNOR2_X1 U6901 ( .A(rs_exe[0]), .B(n7538), .ZN(n5269) );
  XNOR2_X1 U6902 ( .A(rs_exe[1]), .B(n7537), .ZN(n5270) );
  XNOR2_X1 U6903 ( .A(rs_exe[3]), .B(n7535), .ZN(n5267) );
  XNOR2_X1 U6904 ( .A(rs_exe[4]), .B(n7534), .ZN(n5271) );
  XNOR2_X1 U6905 ( .A(rs_exe[2]), .B(n7536), .ZN(n5268) );
  INV_X1 U6906 ( .A(n5340), .ZN(n4835) );
  XNOR2_X1 U6907 ( .A(rs_exe[3]), .B(rd_exemem[3]), .ZN(n5263) );
  NAND3_X1 U6908 ( .A1(n5238), .A2(n4794), .A3(n5237), .ZN(n4744) );
  AND2_X1 U6909 ( .A1(\ctrl_u/curr_exe_40 ), .A2(\ctrl_u/curr_wb[3] ), .ZN(
        n5237) );
  XNOR2_X1 U6910 ( .A(rt_exe[3]), .B(n7535), .ZN(n5238) );
  NAND3_X1 U6911 ( .A1(n5236), .A2(n5235), .A3(n4793), .ZN(n4743) );
  XNOR2_X1 U6912 ( .A(rt_exe[4]), .B(n7534), .ZN(n5235) );
  XNOR2_X1 U6913 ( .A(rt_exe[2]), .B(n7536), .ZN(n5236) );
  AND2_X1 U6914 ( .A1(n7171), .A2(en_imm_id), .ZN(n7151) );
  INV_X1 U6915 ( .A(shift_reg_id), .ZN(n6896) );
  INV_X1 U6916 ( .A(en_rd_id), .ZN(n7140) );
  INV_X1 U6917 ( .A(en_b_id), .ZN(n5011) );
  INV_X1 U6918 ( .A(en_a_neg_id), .ZN(n6334) );
  AND2_X1 U6919 ( .A1(en_shift_reg_id), .A2(n6896), .ZN(n4111) );
  INV_X1 U6920 ( .A(n5215), .ZN(n4682) );
  INV_X1 U6921 ( .A(\ctrl_u/if_stall ), .ZN(n4934) );
  OR2_X1 U6922 ( .A1(\ctrl_u/if_stall ), .A2(n5339), .ZN(n4117) );
  INV_X1 U6923 ( .A(n6416), .ZN(n4899) );
  OR2_X1 U6924 ( .A1(n4356), .A2(n4221), .ZN(n4122) );
  OAI21_X1 U6925 ( .B1(n7260), .B2(n4262), .A(n7257), .ZN(n99) );
  INV_X1 U6926 ( .A(n6449), .ZN(n4887) );
  AND2_X1 U6927 ( .A1(\dp/npc_id_exe_int[4] ), .A2(\dp/imm_id_exe_int[4] ), 
        .ZN(n4129) );
  INV_X1 U6928 ( .A(n7437), .ZN(n4891) );
  INV_X1 U6929 ( .A(n7106), .ZN(n4892) );
  INV_X1 U6930 ( .A(n6447), .ZN(n4888) );
  AND2_X1 U6931 ( .A1(\dp/npc_id_exe_int[25] ), .A2(n4124), .ZN(n4131) );
  NOR2_X1 U6932 ( .A1(\ctrl_u/if_stall ), .A2(n4646), .ZN(n5038) );
  NOR2_X1 U6933 ( .A1(\ctrl_u/curr_id[17] ), .A2(\ctrl_u/n70 ), .ZN(n4132) );
  NOR2_X1 U6934 ( .A1(n3873), .A2(n4356), .ZN(n4133) );
  INV_X1 U6935 ( .A(n6306), .ZN(n6308) );
  AND2_X1 U6936 ( .A1(n4111), .A2(b_selector_id), .ZN(n4134) );
  AND2_X1 U6937 ( .A1(n4111), .A2(n4357), .ZN(n4135) );
  NOR2_X1 U6938 ( .A1(n3915), .A2(n6182), .ZN(n5192) );
  INV_X1 U6939 ( .A(n7258), .ZN(n4715) );
  NAND2_X1 U6940 ( .A1(n5922), .A2(n5921), .ZN(n5091) );
  AOI21_X1 U6941 ( .B1(n5617), .B2(n3924), .A(n7340), .ZN(n5343) );
  INV_X1 U6942 ( .A(n5343), .ZN(n4867) );
  OAI21_X1 U6943 ( .B1(n7260), .B2(n4263), .A(n4715), .ZN(n95) );
  NAND2_X1 U6944 ( .A1(n4037), .A2(n4726), .ZN(n5658) );
  AND2_X1 U6945 ( .A1(\dp/npc_id_exe_int[23] ), .A2(\dp/imm_id_exe_int[23] ), 
        .ZN(n4275) );
  AND2_X1 U6946 ( .A1(\dp/npc_id_exe_int[17] ), .A2(n4115), .ZN(n4276) );
  INV_X1 U6947 ( .A(n5940), .ZN(n4958) );
  INV_X1 U6948 ( .A(n6419), .ZN(n4895) );
  INV_X1 U6949 ( .A(\intadd_1/n56 ), .ZN(n4751) );
  NAND2_X1 U6950 ( .A1(n7171), .A2(en_npc_id), .ZN(n7139) );
  INV_X1 U6951 ( .A(n6417), .ZN(n4901) );
  INV_X1 U6952 ( .A(n6418), .ZN(n4897) );
  INV_X1 U6953 ( .A(n7438), .ZN(n4910) );
  INV_X1 U6954 ( .A(n6434), .ZN(n4890) );
  AOI21_X1 U6955 ( .B1(\dp/exs/alu_unit/shifter_out[3] ), .B2(n7083), .A(n5835), .ZN(n6464) );
  INV_X1 U6956 ( .A(n6464), .ZN(n4881) );
  INV_X1 U6957 ( .A(n6462), .ZN(n4882) );
  AOI21_X1 U6958 ( .B1(\dp/exs/alu_unit/shifter_out[5] ), .B2(n7083), .A(n5863), .ZN(n6460) );
  INV_X1 U6959 ( .A(n6460), .ZN(n4883) );
  INV_X1 U6960 ( .A(n6457), .ZN(n4884) );
  AOI21_X1 U6961 ( .B1(\dp/exs/alu_unit/shifter_out[7] ), .B2(n3954), .A(n5892), .ZN(n6454) );
  INV_X1 U6962 ( .A(n6454), .ZN(n4885) );
  INV_X1 U6963 ( .A(n6451), .ZN(n4886) );
  INV_X1 U6964 ( .A(n6445), .ZN(n4889) );
  AOI21_X1 U6965 ( .B1(n6053), .B2(n7076), .A(n6052), .ZN(n6420) );
  INV_X1 U6966 ( .A(n6420), .ZN(n4893) );
  INV_X1 U6967 ( .A(n6421), .ZN(n4900) );
  INV_X1 U6968 ( .A(pc_en), .ZN(n5422) );
  AND2_X1 U6969 ( .A1(n4208), .A2(\intadd_1/n45 ), .ZN(n4288) );
  OR2_X1 U6970 ( .A1(n6494), .A2(n6493), .ZN(n4289) );
  OR2_X1 U6971 ( .A1(n6592), .A2(n6591), .ZN(n4290) );
  AND2_X1 U6972 ( .A1(\intadd_1/n183 ), .A2(\intadd_1/n83 ), .ZN(n4296) );
  AND3_X1 U6973 ( .A1(\dp/b_mult_id_exe_int[2] ), .A2(n594), .A3(n595), .ZN(
        n4297) );
  INV_X1 U6974 ( .A(n5100), .ZN(n5957) );
  OR2_X1 U6975 ( .A1(n6089), .A2(n6090), .ZN(n4309) );
  OR2_X1 U6976 ( .A1(n5970), .A2(n5971), .ZN(n4310) );
  AND2_X1 U6977 ( .A1(n3936), .A2(\dp/pc_plus4_out_if_int[21] ), .ZN(n4311) );
  AND2_X1 U6978 ( .A1(n3936), .A2(\dp/pc_plus4_out_if_int[23] ), .ZN(n4312) );
  AND2_X1 U6979 ( .A1(n3936), .A2(\dp/pc_plus4_out_if_int[24] ), .ZN(n4313) );
  AND2_X1 U6980 ( .A1(n3928), .A2(\dp/pc_plus4_out_if_int[26] ), .ZN(n4314) );
  NOR2_X1 U6981 ( .A1(n5104), .A2(n5101), .ZN(n5099) );
  OR2_X1 U6982 ( .A1(n6414), .A2(n3885), .ZN(n4315) );
  AND2_X1 U6983 ( .A1(en_b_id), .A2(data_tbs_selector_id), .ZN(n4316) );
  OR2_X1 U6984 ( .A1(\intadd_2/SUM[22] ), .A2(n3937), .ZN(n4319) );
  INV_X1 U6985 ( .A(n6701), .ZN(n5124) );
  NOR2_X1 U6986 ( .A1(\intadd_1/A[28] ), .A2(\intadd_1/B[28] ), .ZN(n4320) );
  AND2_X1 U6987 ( .A1(n5193), .A2(btb_cache_read_address[28]), .ZN(n4321) );
  NAND2_X1 U6988 ( .A1(pc_en), .A2(rst_mem_wb_regs), .ZN(n6181) );
  INV_X1 U6989 ( .A(n6181), .ZN(n6178) );
  AND2_X1 U6990 ( .A1(n5343), .A2(rst_mem_wb_regs), .ZN(n4323) );
  NOR2_X1 U6991 ( .A1(n6004), .A2(n6005), .ZN(n4324) );
  AND2_X1 U6992 ( .A1(\intadd_1/n182 ), .A2(\intadd_1/n78 ), .ZN(n4325) );
  INV_X1 U6993 ( .A(n5020), .ZN(n4999) );
  OR2_X1 U6994 ( .A1(\intadd_2/SUM[23] ), .A2(n3937), .ZN(n4326) );
  OR2_X1 U6995 ( .A1(\intadd_2/SUM[25] ), .A2(n3937), .ZN(n4327) );
  AND2_X1 U6996 ( .A1(n4943), .A2(n5024), .ZN(n4328) );
  OR2_X1 U6997 ( .A1(n6487), .A2(n6488), .ZN(n4329) );
  NAND2_X1 U6998 ( .A1(n5001), .A2(n4796), .ZN(n4331) );
  INV_X1 U6999 ( .A(wp_data[9]), .ZN(n5312) );
  OR2_X1 U7000 ( .A1(n4820), .A2(n6996), .ZN(n4332) );
  OR2_X1 U7001 ( .A1(n4820), .A2(n7001), .ZN(n4333) );
  NAND4_X1 U7002 ( .A1(n6155), .A2(n6154), .A3(n6153), .A4(n6152), .ZN(n6307)
         );
  OR2_X1 U7003 ( .A1(n4820), .A2(n7054), .ZN(n4334) );
  NAND2_X1 U7004 ( .A1(n4835), .A2(n4303), .ZN(n5081) );
  NAND2_X1 U7005 ( .A1(\intadd_1/A[25] ), .A2(\intadd_1/B[25] ), .ZN(
        \intadd_1/n33 ) );
  AND2_X1 U7006 ( .A1(n4225), .A2(n4330), .ZN(n4350) );
  INV_X1 U7007 ( .A(n4787), .ZN(n4786) );
  NAND2_X1 U7008 ( .A1(\dp/npc_id_exe_int[5] ), .A2(n4125), .ZN(n4351) );
  AND2_X1 U7009 ( .A1(en_shift_reg_id), .A2(shift_reg_id), .ZN(n4353) );
  INV_X1 U7010 ( .A(en_mul_id), .ZN(n6721) );
  AND2_X1 U7011 ( .A1(n4943), .A2(n5025), .ZN(n4354) );
  OR2_X1 U7012 ( .A1(n4747), .A2(n4131), .ZN(n4355) );
  NAND2_X1 U7013 ( .A1(n5751), .A2(log_type_exe[1]), .ZN(n6157) );
  XOR2_X1 U7014 ( .A(\dp/npc_id_exe_int[31] ), .B(\dp/imm_id_exe_int[31] ), 
        .Z(n4449) );
  OR2_X1 U7015 ( .A1(n6981), .A2(n4402), .ZN(n4603) );
  NAND3_X1 U7016 ( .A1(instr_if[3]), .A2(n7281), .A3(n5534), .ZN(n4604) );
  NAND2_X1 U7017 ( .A1(n5540), .A2(n5537), .ZN(n4605) );
  NOR3_X1 U7018 ( .A1(instr_if[5]), .A2(n5577), .A3(n7279), .ZN(n5480) );
  OR2_X1 U7019 ( .A1(instr_if[29]), .A2(n5548), .ZN(n4646) );
  AND2_X1 U7020 ( .A1(n5513), .A2(n5605), .ZN(n4647) );
  NAND2_X1 U7021 ( .A1(n6971), .A2(n4684), .ZN(n2728) );
  NAND2_X1 U7022 ( .A1(n6982), .A2(n4685), .ZN(n2732) );
  NAND2_X1 U7023 ( .A1(n6986), .A2(n4686), .ZN(n2735) );
  NAND2_X1 U7024 ( .A1(n6994), .A2(n4687), .ZN(n2738) );
  NAND2_X1 U7025 ( .A1(n6973), .A2(n4688), .ZN(n2729) );
  NAND2_X1 U7026 ( .A1(n6983), .A2(n4689), .ZN(n2733) );
  NAND2_X1 U7027 ( .A1(n6988), .A2(n4690), .ZN(n2736) );
  NAND2_X1 U7028 ( .A1(n6969), .A2(n4691), .ZN(n2727) );
  NAND2_X1 U7029 ( .A1(n6977), .A2(n4692), .ZN(n2730) );
  NAND2_X1 U7030 ( .A1(n6990), .A2(n4694), .ZN(n2737) );
  NAND2_X1 U7031 ( .A1(n7011), .A2(n4695), .ZN(n2742) );
  NAND2_X1 U7032 ( .A1(n6984), .A2(n4693), .ZN(n2734) );
  NAND2_X1 U7033 ( .A1(n4648), .A2(rt_id[3]), .ZN(n4673) );
  AOI21_X1 U7034 ( .B1(n3931), .B2(\dp/ifs/pc_btb[17] ), .A(n4649), .ZN(n6392)
         );
  OAI21_X1 U7035 ( .B1(n3873), .B2(n4110), .A(n4650), .ZN(n4649) );
  NAND2_X1 U7036 ( .A1(n7108), .A2(btb_cache_read_address[17]), .ZN(n4650) );
  AOI21_X1 U7037 ( .B1(n3894), .B2(\dp/ifs/pc_btb[16] ), .A(n4652), .ZN(n6390)
         );
  OAI21_X1 U7038 ( .B1(n3873), .B2(n4113), .A(n4653), .ZN(n4652) );
  NAND2_X1 U7039 ( .A1(n5193), .A2(btb_cache_read_address[16]), .ZN(n4653) );
  AOI21_X1 U7040 ( .B1(n3894), .B2(\dp/ifs/pc_btb[18] ), .A(n4654), .ZN(n6394)
         );
  OAI21_X1 U7041 ( .B1(n3873), .B2(n4114), .A(n4655), .ZN(n4654) );
  NAND2_X1 U7042 ( .A1(n5193), .A2(btb_cache_read_address[18]), .ZN(n4655) );
  AOI21_X1 U7043 ( .B1(n3894), .B2(\dp/ifs/pc_btb[10] ), .A(n4656), .ZN(n6373)
         );
  OAI21_X1 U7044 ( .B1(n3873), .B2(n4234), .A(n4657), .ZN(n4656) );
  NAND2_X1 U7045 ( .A1(n7108), .A2(btb_cache_read_address[10]), .ZN(n4657) );
  OAI21_X1 U7046 ( .B1(n5565), .B2(\ctrl_u/curr_id[14] ), .A(n5564), .ZN(
        \ctrl_u/n384 ) );
  OAI21_X1 U7047 ( .B1(n5565), .B2(\ctrl_u/curr_id[5] ), .A(n5564), .ZN(
        \ctrl_u/n406 ) );
  OAI21_X1 U7048 ( .B1(n5565), .B2(\ctrl_u/curr_id[1] ), .A(n5564), .ZN(
        \ctrl_u/n412 ) );
  AOI21_X1 U7049 ( .B1(n3895), .B2(\dp/ifs/pc_btb[11] ), .A(n4658), .ZN(n6375)
         );
  OAI21_X1 U7050 ( .B1(n3873), .B2(n4226), .A(n4659), .ZN(n4658) );
  NAND2_X1 U7051 ( .A1(n7108), .A2(btb_cache_read_address[11]), .ZN(n4659) );
  NAND2_X1 U7052 ( .A1(n4315), .A2(n4660), .ZN(n2530) );
  NOR2_X1 U7053 ( .A1(n4663), .A2(n4661), .ZN(n4660) );
  INV_X1 U7054 ( .A(\intadd_2/SUM[26] ), .ZN(n4662) );
  INV_X1 U7055 ( .A(n6404), .ZN(n4663) );
  AOI21_X1 U7056 ( .B1(n3895), .B2(\dp/ifs/pc_btb[12] ), .A(n4665), .ZN(n6377)
         );
  OAI21_X1 U7057 ( .B1(n3873), .B2(n4235), .A(n4666), .ZN(n4665) );
  NAND2_X1 U7058 ( .A1(n5193), .A2(btb_cache_read_address[12]), .ZN(n4666) );
  NAND2_X1 U7059 ( .A1(n4667), .A2(n4815), .ZN(\ctrl_u/n528 ) );
  OAI21_X1 U7060 ( .B1(\intadd_1/n159 ), .B2(\intadd_1/n153 ), .A(
        \intadd_1/n154 ), .ZN(\intadd_1/n152 ) );
  AOI21_X1 U7061 ( .B1(n4285), .B2(n5325), .A(n7241), .ZN(\intadd_1/B[4] ) );
  NAND2_X1 U7062 ( .A1(n5122), .A2(n4350), .ZN(n4669) );
  NAND2_X1 U7063 ( .A1(n5260), .A2(n4225), .ZN(n4670) );
  OR2_X1 U7064 ( .A1(n5260), .A2(n4225), .ZN(n4671) );
  XNOR2_X1 U7065 ( .A(n5144), .B(n4225), .ZN(\intadd_1/A[8] ) );
  NAND4_X1 U7066 ( .A1(n6914), .A2(n6958), .A3(n6915), .A4(n4673), .ZN(n2698)
         );
  NAND2_X1 U7067 ( .A1(n4674), .A2(n4815), .ZN(\ctrl_u/n527 ) );
  NAND2_X1 U7068 ( .A1(n3932), .A2(n4135), .ZN(n6947) );
  OAI22_X1 U7069 ( .A1(n4071), .A2(n5173), .B1(n5172), .B2(n5319), .ZN(n7243)
         );
  XNOR2_X1 U7070 ( .A(n6036), .B(sub_add_exe), .ZN(n4699) );
  XNOR2_X1 U7071 ( .A(n5995), .B(sub_add_exe), .ZN(\intadd_1/A[19] ) );
  AOI21_X1 U7072 ( .B1(n5135), .B2(n4337), .A(n4701), .ZN(n5995) );
  OAI22_X1 U7073 ( .A1(n3913), .A2(wp_data[20]), .B1(
        \dp/mul_feedback_exe_mem_int[20] ), .B2(n3922), .ZN(n4701) );
  XNOR2_X1 U7074 ( .A(n6012), .B(sub_add_exe), .ZN(n4845) );
  OAI22_X1 U7075 ( .A1(n4040), .A2(wp_data[21]), .B1(n3922), .B2(
        \dp/mul_feedback_exe_mem_int[21] ), .ZN(n4702) );
  NAND3_X1 U7076 ( .A1(n4266), .A2(cpu_is_reading), .A3(\ctrl_u/curr_ms ), 
        .ZN(n4704) );
  INV_X1 U7077 ( .A(n5119), .ZN(n4705) );
  NAND2_X1 U7078 ( .A1(n5308), .A2(n5307), .ZN(n7229) );
  NAND2_X1 U7079 ( .A1(n4708), .A2(n4788), .ZN(n4707) );
  NAND2_X1 U7080 ( .A1(\intadd_1/n30 ), .A2(n4803), .ZN(n4708) );
  NAND2_X1 U7081 ( .A1(n4732), .A2(n4775), .ZN(\intadd_1/n30 ) );
  XNOR2_X1 U7082 ( .A(n4761), .B(n4325), .ZN(\intadd_1/SUM[17] ) );
  XNOR2_X1 U7083 ( .A(\intadd_1/n46 ), .B(n4288), .ZN(\intadd_1/SUM[23] ) );
  XNOR2_X1 U7084 ( .A(rs_exe[2]), .B(rd_exemem[2]), .ZN(n4710) );
  XNOR2_X1 U7085 ( .A(rs_exe[4]), .B(rd_exemem[4]), .ZN(n4711) );
  OAI211_X1 U7086 ( .C1(n4714), .C2(n4733), .A(n4713), .B(n4712), .ZN(
        \intadd_1/A[0] ) );
  NAND2_X1 U7087 ( .A1(n7258), .A2(sub_add_exe), .ZN(n4712) );
  NAND2_X1 U7088 ( .A1(n4733), .A2(sub_add_exe), .ZN(n4713) );
  OR2_X1 U7089 ( .A1(n7258), .A2(sub_add_exe), .ZN(n4714) );
  NAND2_X1 U7090 ( .A1(n6089), .A2(n6090), .ZN(n4716) );
  NAND2_X1 U7091 ( .A1(n6088), .A2(n4309), .ZN(n4717) );
  NAND2_X1 U7092 ( .A1(n4719), .A2(n4718), .ZN(n6088) );
  NAND2_X1 U7093 ( .A1(n6075), .A2(n6074), .ZN(n4718) );
  OAI21_X1 U7094 ( .B1(n6075), .B2(n6074), .A(n6073), .ZN(n4719) );
  INV_X1 U7095 ( .A(n4720), .ZN(\intadd_1/n131 ) );
  NAND2_X1 U7096 ( .A1(n4229), .A2(\intadd_1/n37 ), .ZN(n4724) );
  INV_X1 U7097 ( .A(\intadd_1/n39 ), .ZN(n4725) );
  NAND3_X1 U7098 ( .A1(n4726), .A2(n4037), .A3(n4232), .ZN(n5142) );
  NAND4_X1 U7099 ( .A1(n3961), .A2(n4726), .A3(n4037), .A4(n5097), .ZN(n5171)
         );
  NAND2_X1 U7100 ( .A1(\intadd_1/SUM[27] ), .A2(\intadd_1/SUM[21] ), .ZN(n4770) );
  XNOR2_X1 U7101 ( .A(n4727), .B(n4298), .ZN(\intadd_1/SUM[21] ) );
  OAI21_X1 U7102 ( .B1(n4760), .B2(n4759), .A(n4756), .ZN(n4727) );
  XNOR2_X1 U7103 ( .A(\intadd_1/n30 ), .B(n4804), .ZN(\intadd_1/SUM[27] ) );
  XNOR2_X1 U7104 ( .A(\intadd_1/n84 ), .B(n4296), .ZN(\intadd_1/SUM[16] ) );
  AND2_X1 U7105 ( .A1(n4959), .A2(n4303), .ZN(n4735) );
  XNOR2_X1 U7106 ( .A(rt_exe[2]), .B(rd_exemem[2]), .ZN(n4842) );
  NAND2_X1 U7107 ( .A1(n5063), .A2(n5088), .ZN(n4741) );
  OAI21_X1 U7108 ( .B1(n3957), .B2(n4355), .A(n4745), .ZN(\intadd_2/n6 ) );
  XNOR2_X1 U7109 ( .A(n4749), .B(n4748), .ZN(\intadd_2/SUM[22] ) );
  INV_X1 U7110 ( .A(\intadd_1/n60 ), .ZN(n4757) );
  INV_X1 U7111 ( .A(\intadd_1/n59 ), .ZN(n4758) );
  NAND2_X1 U7112 ( .A1(\intadd_1/n68 ), .A2(n3863), .ZN(n4759) );
  XNOR2_X1 U7113 ( .A(\intadd_1/n55 ), .B(\intadd_1/n4 ), .ZN(
        \intadd_1/SUM[22] ) );
  NAND2_X1 U7114 ( .A1(n4782), .A2(n4780), .ZN(n5969) );
  INV_X1 U7115 ( .A(n4781), .ZN(n4780) );
  NOR2_X1 U7116 ( .A1(n5099), .A2(n4785), .ZN(n4783) );
  NAND2_X1 U7117 ( .A1(n5943), .A2(n5942), .ZN(n4787) );
  NAND2_X1 U7118 ( .A1(n4792), .A2(n5340), .ZN(n5086) );
  NOR2_X1 U7119 ( .A1(n4837), .A2(n4838), .ZN(n4792) );
  XNOR2_X1 U7120 ( .A(rt_exe[1]), .B(n7537), .ZN(n4793) );
  XNOR2_X1 U7121 ( .A(n3904), .B(n7538), .ZN(n4794) );
  NAND2_X1 U7122 ( .A1(n5182), .A2(n5549), .ZN(n5564) );
  NAND2_X1 U7123 ( .A1(n3902), .A2(n5011), .ZN(n6931) );
  INV_X1 U7124 ( .A(n3929), .ZN(n5619) );
  AOI21_X1 U7125 ( .B1(n4832), .B2(\intadd_1/n107 ), .A(\intadd_1/n108 ), .ZN(
        n4831) );
  INV_X1 U7126 ( .A(\intadd_1/n119 ), .ZN(n4832) );
  NAND2_X1 U7127 ( .A1(n4834), .A2(\intadd_1/n107 ), .ZN(n4833) );
  INV_X1 U7128 ( .A(\intadd_1/n118 ), .ZN(n4834) );
  NAND4_X1 U7129 ( .A1(n5268), .A2(n5271), .A3(n5267), .A4(\ctrl_u/curr_wb[3] ), .ZN(n4837) );
  NAND2_X1 U7130 ( .A1(n5270), .A2(n5269), .ZN(n4838) );
  INV_X1 U7131 ( .A(en_add_id), .ZN(n4843) );
  NOR2_X1 U7132 ( .A1(n4052), .A2(n4851), .ZN(n5510) );
  NAND2_X1 U7133 ( .A1(n4853), .A2(n4852), .ZN(n4851) );
  AOI21_X1 U7134 ( .B1(n3859), .B2(n4117), .A(n4647), .ZN(n4852) );
  NAND2_X1 U7135 ( .A1(n4854), .A2(n4117), .ZN(n4853) );
  INV_X1 U7136 ( .A(en_shift_reg_id), .ZN(n4855) );
  NAND3_X1 U7137 ( .A1(n4933), .A2(n4850), .A3(n5481), .ZN(n5488) );
  NOR2_X1 U7138 ( .A1(n6182), .A2(n6181), .ZN(n4875) );
  NOR2_X1 U7139 ( .A1(n4878), .A2(n4877), .ZN(n6399) );
  NOR2_X1 U7140 ( .A1(n3873), .A2(n4103), .ZN(n4878) );
  OAI211_X1 U7141 ( .C1(n4988), .C2(\intadd_1/n28 ), .A(n4880), .B(n4961), 
        .ZN(n6164) );
  NAND2_X1 U7142 ( .A1(\intadd_1/n28 ), .A2(n4987), .ZN(n4880) );
  INV_X1 U7143 ( .A(n4907), .ZN(n4906) );
  OAI21_X1 U7144 ( .B1(\intadd_1/n28 ), .B2(n4983), .A(n5335), .ZN(n4907) );
  XNOR2_X1 U7145 ( .A(n4912), .B(n4289), .ZN(n6495) );
  XNOR2_X1 U7146 ( .A(n4915), .B(n4290), .ZN(n6593) );
  OAI21_X1 U7147 ( .B1(n6701), .B2(n4917), .A(n4916), .ZN(n4915) );
  AOI21_X1 U7148 ( .B1(n6588), .B2(n6589), .A(n6587), .ZN(n4916) );
  NAND2_X1 U7149 ( .A1(n6586), .A2(n6589), .ZN(n4917) );
  AOI21_X1 U7150 ( .B1(\intadd_2/n17 ), .B2(n4926), .A(n4924), .ZN(n4923) );
  NAND2_X1 U7151 ( .A1(n4940), .A2(n4939), .ZN(n4938) );
  NAND2_X1 U7152 ( .A1(n5119), .A2(n4344), .ZN(n4939) );
  INV_X1 U7153 ( .A(n5251), .ZN(n4940) );
  NAND2_X1 U7154 ( .A1(\dp/npc_id_exe_int[21] ), .A2(\dp/imm_id_exe_int[21] ), 
        .ZN(n4941) );
  INV_X1 U7155 ( .A(n7092), .ZN(n4945) );
  NOR2_X1 U7156 ( .A1(n4955), .A2(n4952), .ZN(n4950) );
  XNOR2_X1 U7157 ( .A(rt_exe[4]), .B(rd_exemem[4]), .ZN(n4959) );
  NAND2_X1 U7158 ( .A1(n6406), .A2(n4963), .ZN(n4962) );
  AOI21_X1 U7159 ( .B1(n3895), .B2(\dp/ifs/pc_btb[28] ), .A(n4321), .ZN(n4963)
         );
  NAND2_X1 U7160 ( .A1(n4969), .A2(n4319), .ZN(n2534) );
  AOI211_X1 U7161 ( .C1(n6405), .C2(\dp/npc_id_exe_int[25] ), .A(n4970), .B(
        n4312), .ZN(n4969) );
  AOI21_X1 U7162 ( .B1(n4054), .B2(\dp/ifs/pc_btb[23] ), .A(n4972), .ZN(n4971)
         );
  NOR2_X1 U7163 ( .A1(n6402), .A2(n4596), .ZN(n4972) );
  NAND2_X1 U7164 ( .A1(n4326), .A2(n4973), .ZN(n2533) );
  AOI211_X1 U7165 ( .C1(n6405), .C2(\dp/npc_id_exe_int[26] ), .A(n4974), .B(
        n4313), .ZN(n4973) );
  AOI21_X1 U7166 ( .B1(n4054), .B2(\dp/ifs/pc_btb[24] ), .A(n4976), .ZN(n4975)
         );
  NOR2_X1 U7167 ( .A1(n6402), .A2(n4597), .ZN(n4976) );
  NAND2_X1 U7168 ( .A1(n4327), .A2(n4977), .ZN(n2531) );
  AOI211_X1 U7169 ( .C1(n6405), .C2(\dp/npc_id_exe_int[28] ), .A(n4314), .B(
        n4978), .ZN(n4977) );
  AOI21_X1 U7170 ( .B1(n4054), .B2(\dp/ifs/pc_btb[26] ), .A(n4980), .ZN(n4979)
         );
  NOR2_X1 U7171 ( .A1(n6402), .A2(n4598), .ZN(n4980) );
  NAND2_X1 U7172 ( .A1(\intadd_1/n28 ), .A2(n4982), .ZN(n4981) );
  OAI21_X1 U7173 ( .B1(n4986), .B2(n4987), .A(n5071), .ZN(n4982) );
  INV_X1 U7174 ( .A(n4984), .ZN(n4983) );
  OAI21_X1 U7175 ( .B1(n4986), .B2(n5049), .A(n4985), .ZN(n4984) );
  INV_X1 U7176 ( .A(n5071), .ZN(n4985) );
  NAND2_X1 U7177 ( .A1(n5928), .A2(n5929), .ZN(n4990) );
  OR2_X1 U7178 ( .A1(n5928), .A2(n5929), .ZN(n4991) );
  OAI21_X1 U7179 ( .B1(n4998), .B2(n4017), .A(n4996), .ZN(\intadd_2/n23 ) );
  INV_X1 U7180 ( .A(n4997), .ZN(n4996) );
  OAI21_X1 U7181 ( .B1(n5039), .B2(n4999), .A(n5019), .ZN(n4997) );
  NAND2_X1 U7182 ( .A1(n5040), .A2(n5020), .ZN(n4998) );
  NAND2_X1 U7183 ( .A1(n4116), .A2(\dp/imm_id_exe_int[15] ), .ZN(n5002) );
  INV_X1 U7184 ( .A(n6184), .ZN(n5009) );
  XNOR2_X1 U7185 ( .A(n5010), .B(n4449), .ZN(n5087) );
  AOI22_X1 U7186 ( .A1(\intadd_2/n2 ), .A2(n5013), .B1(n4367), .B2(n4519), 
        .ZN(n5010) );
  NAND2_X1 U7187 ( .A1(n4140), .A2(\dp/imm_id_exe_int[30] ), .ZN(n5013) );
  NAND2_X1 U7188 ( .A1(n4216), .A2(n4098), .ZN(n5019) );
  NAND2_X1 U7189 ( .A1(\dp/npc_id_exe_int[8] ), .A2(\dp/imm_id_exe_int[8] ), 
        .ZN(n5020) );
  INV_X1 U7190 ( .A(n5064), .ZN(n5032) );
  NAND3_X1 U7191 ( .A1(n5046), .A2(n5045), .A3(\ctrl_u/curr_exe[19] ), .ZN(
        n6177) );
  NAND2_X1 U7192 ( .A1(n4123), .A2(cond_sel_exe[1]), .ZN(n5042) );
  NOR2_X1 U7193 ( .A1(n4123), .A2(cond_sel_exe[1]), .ZN(n5043) );
  NAND2_X1 U7194 ( .A1(n5821), .A2(btb_cache_update_data), .ZN(n5046) );
  NOR2_X1 U7195 ( .A1(n6402), .A2(n4599), .ZN(n5047) );
  OAI211_X1 U7196 ( .C1(n5084), .C2(n5057), .A(n4351), .B(n5055), .ZN(n5054)
         );
  NAND2_X1 U7197 ( .A1(n4129), .A2(n5082), .ZN(n5055) );
  NAND2_X1 U7198 ( .A1(n5058), .A2(\intadd_1/n65 ), .ZN(\intadd_1/n63 ) );
  INV_X1 U7199 ( .A(\intadd_1/n64 ), .ZN(n5059) );
  INV_X1 U7200 ( .A(n5070), .ZN(n5069) );
  OAI211_X1 U7201 ( .C1(\intadd_2/SUM[27] ), .C2(n6167), .A(n6132), .B(n6131), 
        .ZN(btb_cache_data_in[28]) );
  NAND2_X1 U7202 ( .A1(n4215), .A2(n4099), .ZN(n5072) );
  NAND2_X1 U7203 ( .A1(\dp/npc_id_exe_int[6] ), .A2(\dp/imm_id_exe_int[6] ), 
        .ZN(n5073) );
  NAND2_X1 U7204 ( .A1(n4209), .A2(\intadd_2/A[2] ), .ZN(n5078) );
  NAND2_X1 U7205 ( .A1(n5085), .A2(n5093), .ZN(n5084) );
  NAND2_X1 U7206 ( .A1(n4214), .A2(n4100), .ZN(n5082) );
  OAI21_X1 U7207 ( .B1(n4213), .B2(\intadd_2/A[0] ), .A(n5095), .ZN(n5085) );
  NAND2_X1 U7208 ( .A1(\dp/npc_id_exe_int[2] ), .A2(\dp/imm_id_exe_int[2] ), 
        .ZN(n5095) );
  INV_X1 U7209 ( .A(n5091), .ZN(n5089) );
  NAND2_X1 U7210 ( .A1(n4213), .A2(\intadd_2/A[0] ), .ZN(n5093) );
  NOR3_X1 U7212 ( .A1(n4031), .A2(n5767), .A3(n4300), .ZN(op_b_fw_sel_exe[1])
         );
  NAND2_X1 U7213 ( .A1(\intadd_1/A[5] ), .A2(\intadd_1/B[5] ), .ZN(
        \intadd_1/n149 ) );
  NAND2_X1 U7214 ( .A1(\intadd_1/A[19] ), .A2(\intadd_1/B[19] ), .ZN(
        \intadd_1/n65 ) );
  NOR3_X1 U7215 ( .A1(n7188), .A2(n5229), .A3(\mc/currstate[0] ), .ZN(n3114)
         );
  XNOR2_X1 U7216 ( .A(n5752), .B(n4225), .ZN(\intadd_1/A[15] ) );
  NOR2_X1 U7217 ( .A1(n7065), .A2(n7064), .ZN(n7070) );
  OR2_X1 U7218 ( .A1(n7064), .A2(n7071), .ZN(n7079) );
  NOR2_X1 U7219 ( .A1(n7253), .A2(n463), .ZN(n5327) );
  NAND2_X1 U7220 ( .A1(\intadd_1/n143 ), .A2(\intadd_1/n151 ), .ZN(
        \intadd_1/n141 ) );
  NAND2_X1 U7221 ( .A1(\intadd_1/A[2] ), .A2(\intadd_1/B[2] ), .ZN(
        \intadd_1/n165 ) );
  AOI22_X1 U7222 ( .A1(n6413), .A2(n5194), .B1(\dp/a_neg_mult_id_exe_int[30] ), 
        .B2(n5126), .ZN(n1446) );
  NAND2_X1 U7223 ( .A1(n6413), .A2(n3884), .ZN(n6407) );
  OAI21_X1 U7224 ( .B1(n6701), .B2(n6548), .A(n6547), .ZN(n6544) );
  OAI21_X1 U7225 ( .B1(n6701), .B2(n6684), .A(n6683), .ZN(n6688) );
  OAI22_X1 U7226 ( .A1(n6604), .A2(n7062), .B1(n4193), .B2(n3938), .ZN(n2801)
         );
  OAI22_X1 U7227 ( .A1(n6604), .A2(n5196), .B1(n4488), .B2(n5199), .ZN(n2833)
         );
  OAI22_X1 U7228 ( .A1(n6528), .A2(n7062), .B1(n4189), .B2(n3938), .ZN(n2811)
         );
  OAI22_X1 U7229 ( .A1(n6540), .A2(n7062), .B1(n4190), .B2(n3938), .ZN(n2809)
         );
  OAI22_X1 U7230 ( .A1(n6540), .A2(n5198), .B1(n4504), .B2(n5199), .ZN(n2841)
         );
  OAI22_X1 U7231 ( .A1(n6720), .A2(n7062), .B1(n7435), .B2(n3938), .ZN(n2788)
         );
  OAI22_X1 U7232 ( .A1(n6720), .A2(n5196), .B1(n4585), .B2(n5199), .ZN(n2820)
         );
  OAI22_X1 U7233 ( .A1(n6611), .A2(n7062), .B1(n7433), .B2(n3942), .ZN(n2800)
         );
  OAI22_X1 U7234 ( .A1(n6611), .A2(n5196), .B1(n4407), .B2(n5199), .ZN(n2832)
         );
  OAI22_X1 U7235 ( .A1(n6585), .A2(n7062), .B1(n7432), .B2(n3938), .ZN(n2804)
         );
  OAI22_X1 U7236 ( .A1(n6585), .A2(n5196), .B1(n4486), .B2(n5199), .ZN(n2836)
         );
  OAI22_X1 U7237 ( .A1(n6531), .A2(n7062), .B1(n7431), .B2(n3942), .ZN(n2810)
         );
  OAI22_X1 U7238 ( .A1(n6531), .A2(n5198), .B1(n4505), .B2(n5199), .ZN(n2842)
         );
  OAI22_X1 U7239 ( .A1(n6485), .A2(n7062), .B1(n7430), .B2(n3938), .ZN(n2816)
         );
  OAI22_X1 U7240 ( .A1(n6485), .A2(n5197), .B1(n4480), .B2(n5199), .ZN(n2848)
         );
  OAI22_X1 U7241 ( .A1(n6649), .A2(n7062), .B1(n4195), .B2(n7439), .ZN(n2796)
         );
  XNOR2_X1 U7242 ( .A(n6648), .B(n6647), .ZN(n6649) );
  XNOR2_X1 U7243 ( .A(n6718), .B(n6717), .ZN(n6720) );
  XNOR2_X1 U7244 ( .A(n6610), .B(n6609), .ZN(n6611) );
  XNOR2_X1 U7245 ( .A(n6584), .B(n6583), .ZN(n6585) );
  XNOR2_X1 U7246 ( .A(n6484), .B(n6483), .ZN(n6485) );
  XNOR2_X1 U7247 ( .A(n6530), .B(n6529), .ZN(n6531) );
  OAI22_X1 U7248 ( .A1(n6596), .A2(n7062), .B1(n4192), .B2(n3942), .ZN(n2802)
         );
  XNOR2_X1 U7249 ( .A(n6595), .B(n6594), .ZN(n6596) );
  AOI21_X1 U7250 ( .B1(n6130), .B2(n7076), .A(n6129), .ZN(n6412) );
  AOI211_X1 U7251 ( .C1(n6504), .C2(n6514), .A(n6503), .B(n6502), .ZN(n6508)
         );
  NOR3_X1 U7252 ( .A1(n3886), .A2(n6501), .A3(n6510), .ZN(n6502) );
  AOI211_X1 U7253 ( .C1(n6321), .C2(n6712), .A(n6715), .B(n6320), .ZN(n6332)
         );
  NOR3_X1 U7254 ( .A1(n3872), .A2(n6716), .A3(n6711), .ZN(n6320) );
  AOI211_X1 U7255 ( .C1(n6654), .C2(n6665), .A(n6653), .B(n6652), .ZN(n6659)
         );
  NOR3_X1 U7256 ( .A1(n3872), .A2(n6651), .A3(n6650), .ZN(n6652) );
  AOI211_X1 U7257 ( .C1(n6675), .C2(n6674), .A(n6673), .B(n6672), .ZN(n6680)
         );
  NOR3_X1 U7258 ( .A1(n3872), .A2(n6671), .A3(n6670), .ZN(n6672) );
  AOI211_X1 U7259 ( .C1(n6635), .C2(n6634), .A(n6633), .B(n6632), .ZN(n6640)
         );
  NOR3_X1 U7260 ( .A1(n3886), .A2(n6631), .A3(n6630), .ZN(n6632) );
  AOI211_X1 U7261 ( .C1(n6571), .C2(n6570), .A(n6569), .B(n6568), .ZN(n6576)
         );
  NOR3_X1 U7262 ( .A1(n5125), .A2(n6567), .A3(n6578), .ZN(n6568) );
  AOI211_X1 U7263 ( .C1(n6553), .C2(n6552), .A(n6551), .B(n6550), .ZN(n6558)
         );
  NOR3_X1 U7264 ( .A1(n5125), .A2(n6549), .A3(n6548), .ZN(n6550) );
  AOI211_X1 U7265 ( .C1(n6705), .C2(n6704), .A(n6703), .B(n6702), .ZN(n6709)
         );
  NOR3_X1 U7266 ( .A1(n5125), .A2(n6700), .A3(n6699), .ZN(n6702) );
  OAI22_X1 U7267 ( .A1(n6694), .A2(n5197), .B1(n4537), .B2(n5199), .ZN(n2823)
         );
  OAI22_X1 U7268 ( .A1(n6482), .A2(n7062), .B1(n4188), .B2(n3938), .ZN(n2817)
         );
  AOI211_X1 U7269 ( .C1(n6602), .C2(n6625), .A(n6601), .B(n6600), .ZN(n6603)
         );
  AOI211_X1 U7270 ( .C1(n6526), .C2(n6525), .A(n6524), .B(n6523), .ZN(n6527)
         );
  AOI211_X1 U7271 ( .C1(n6538), .C2(n6563), .A(n6537), .B(n6536), .ZN(n6539)
         );
  OAI211_X1 U7272 ( .C1(n6123), .C2(n6122), .A(n6121), .B(n6120), .ZN(n6130)
         );
  OAI211_X1 U7273 ( .C1(n6133), .C2(n6116), .A(n6115), .B(n6122), .ZN(n6121)
         );
  XNOR2_X1 U7274 ( .A(n5125), .B(n6475), .ZN(n6476) );
  OAI21_X1 U7275 ( .B1(n6701), .B2(n6510), .A(n6496), .ZN(n6499) );
  OAI22_X1 U7276 ( .A1(n5317), .A2(n5171), .B1(n5173), .B2(n6456), .ZN(n7239)
         );
  OR2_X1 U7277 ( .A1(n5171), .A2(n5306), .ZN(n5307) );
  OR2_X1 U7278 ( .A1(n5171), .A2(n5278), .ZN(n5279) );
  OR2_X1 U7279 ( .A1(n5171), .A2(n5295), .ZN(n5296) );
  AOI21_X1 U7280 ( .B1(\intadd_1/n160 ), .B2(\intadd_1/n151 ), .A(
        \intadd_1/n152 ), .ZN(\intadd_1/n150 ) );
  OAI22_X1 U7281 ( .A1(n5305), .A2(n5172), .B1(n5123), .B2(n4088), .ZN(n7227)
         );
  OAI22_X1 U7282 ( .A1(n5294), .A2(n5171), .B1(n5123), .B2(n4085), .ZN(n7215)
         );
  OAI22_X1 U7283 ( .A1(n5291), .A2(n5171), .B1(n5123), .B2(n4086), .ZN(n7209)
         );
  OAI22_X1 U7284 ( .A1(n4084), .A2(n5123), .B1(n5171), .B2(n5288), .ZN(n7203)
         );
  NAND2_X1 U7285 ( .A1(\intadd_1/A[17] ), .A2(\intadd_1/B[17] ), .ZN(
        \intadd_1/n78 ) );
  XNOR2_X1 U7286 ( .A(n5961), .B(sub_add_exe), .ZN(\intadd_1/A[17] ) );
  NAND2_X1 U7287 ( .A1(\intadd_1/n192 ), .A2(\intadd_1/n138 ), .ZN(
        \intadd_1/n19 ) );
  NAND2_X1 U7288 ( .A1(\intadd_1/A[3] ), .A2(\intadd_1/B[3] ), .ZN(
        \intadd_1/n159 ) );
  XNOR2_X1 U7289 ( .A(n5837), .B(n4225), .ZN(\intadd_1/A[3] ) );
  NAND2_X1 U7290 ( .A1(\intadd_1/A[13] ), .A2(\intadd_1/B[13] ), .ZN(
        \intadd_1/n103 ) );
  NAND2_X1 U7291 ( .A1(n5119), .A2(\dp/b_adder_id_exe_int[0] ), .ZN(n5326) );
  NAND2_X1 U7292 ( .A1(\intadd_1/n190 ), .A2(\intadd_1/n128 ), .ZN(
        \intadd_1/n17 ) );
  NAND2_X1 U7293 ( .A1(\intadd_1/A[9] ), .A2(\intadd_1/B[9] ), .ZN(
        \intadd_1/n128 ) );
  XNOR2_X1 U7294 ( .A(\intadd_1/n26 ), .B(\intadd_1/CI ), .ZN(
        \intadd_1/SUM[0] ) );
  NAND2_X1 U7295 ( .A1(n6413), .A2(n6165), .ZN(n6132) );
  AOI22_X1 U7296 ( .A1(n6410), .A2(n6165), .B1(btb_cache_update_data), .B2(
        btb_cache_data_out_rw[29]), .ZN(n6166) );
  OAI21_X1 U7297 ( .B1(n7106), .B2(n5117), .A(n5827), .ZN(btb_cache_data_in[0]) );
  OAI222_X1 U7298 ( .A1(n6112), .A2(n6168), .B1(n5117), .B2(n6416), .C1(n3870), 
        .C2(\intadd_2/SUM[25] ), .ZN(btb_cache_data_in[26]) );
  OAI222_X1 U7299 ( .A1(n6097), .A2(n6168), .B1(n5117), .B2(n6417), .C1(n6167), 
        .C2(\intadd_2/SUM[24] ), .ZN(btb_cache_data_in[25]) );
  OAI222_X1 U7300 ( .A1(n6087), .A2(n6168), .B1(n5117), .B2(n6418), .C1(n3870), 
        .C2(\intadd_2/SUM[23] ), .ZN(btb_cache_data_in[24]) );
  OAI222_X1 U7301 ( .A1(n6072), .A2(n6168), .B1(n5117), .B2(n6419), .C1(n6167), 
        .C2(\intadd_2/SUM[22] ), .ZN(btb_cache_data_in[23]) );
  OAI222_X1 U7302 ( .A1(n6054), .A2(n6168), .B1(n5117), .B2(n6420), .C1(n3870), 
        .C2(\intadd_2/SUM[21] ), .ZN(btb_cache_data_in[22]) );
  OAI222_X1 U7303 ( .A1(n6038), .A2(n6168), .B1(n5117), .B2(n6421), .C1(n6167), 
        .C2(\intadd_2/SUM[20] ), .ZN(btb_cache_data_in[21]) );
  OAI222_X1 U7304 ( .A1(n6028), .A2(n6168), .B1(n5117), .B2(n6422), .C1(n3870), 
        .C2(\intadd_2/SUM[19] ), .ZN(btb_cache_data_in[20]) );
  OAI222_X1 U7305 ( .A1(n6019), .A2(n6168), .B1(n5117), .B2(n6424), .C1(n6167), 
        .C2(\intadd_2/SUM[18] ), .ZN(btb_cache_data_in[19]) );
  OAI222_X1 U7306 ( .A1(n6002), .A2(n6168), .B1(n5117), .B2(n6426), .C1(n3870), 
        .C2(\intadd_2/SUM[17] ), .ZN(btb_cache_data_in[18]) );
  OAI222_X1 U7307 ( .A1(n5985), .A2(n6168), .B1(n5117), .B2(n6428), .C1(n6167), 
        .C2(\intadd_2/SUM[16] ), .ZN(btb_cache_data_in[17]) );
  OAI222_X1 U7308 ( .A1(n5968), .A2(n6168), .B1(n5117), .B2(n6430), .C1(n3870), 
        .C2(\intadd_2/SUM[15] ), .ZN(btb_cache_data_in[16]) );
  OAI222_X1 U7309 ( .A1(n5954), .A2(n6168), .B1(n5117), .B2(n7438), .C1(n6167), 
        .C2(\intadd_2/SUM[14] ), .ZN(btb_cache_data_in[15]) );
  OAI222_X1 U7310 ( .A1(n5953), .A2(n6168), .B1(n5117), .B2(n7437), .C1(n3870), 
        .C2(\intadd_2/SUM[13] ), .ZN(btb_cache_data_in[14]) );
  OAI222_X1 U7311 ( .A1(n5952), .A2(n6168), .B1(n5117), .B2(n6434), .C1(n6167), 
        .C2(\intadd_2/SUM[12] ), .ZN(btb_cache_data_in[13]) );
  OAI222_X1 U7312 ( .A1(n5941), .A2(n6168), .B1(n5117), .B2(n6436), .C1(n3870), 
        .C2(\intadd_2/SUM[11] ), .ZN(btb_cache_data_in[12]) );
  OAI222_X1 U7313 ( .A1(n5938), .A2(n6168), .B1(n5117), .B2(n6439), .C1(n6167), 
        .C2(\intadd_2/SUM[10] ), .ZN(btb_cache_data_in[11]) );
  OAI222_X1 U7314 ( .A1(n5927), .A2(n6168), .B1(n5117), .B2(n6442), .C1(n3870), 
        .C2(\intadd_2/SUM[9] ), .ZN(btb_cache_data_in[10]) );
  OAI222_X1 U7315 ( .A1(n5924), .A2(n6168), .B1(n5117), .B2(n6445), .C1(n6167), 
        .C2(\intadd_2/SUM[8] ), .ZN(btb_cache_data_in[9]) );
  OAI222_X1 U7316 ( .A1(n5920), .A2(n6168), .B1(n5117), .B2(n6447), .C1(n3870), 
        .C2(\intadd_2/SUM[7] ), .ZN(btb_cache_data_in[8]) );
  OAI222_X1 U7317 ( .A1(n5916), .A2(n6168), .B1(n5117), .B2(n6449), .C1(n6167), 
        .C2(\intadd_2/SUM[6] ), .ZN(btb_cache_data_in[7]) );
  OAI222_X1 U7318 ( .A1(n5905), .A2(n6168), .B1(n5117), .B2(n6451), .C1(n3870), 
        .C2(\intadd_2/SUM[5] ), .ZN(btb_cache_data_in[6]) );
  OAI222_X1 U7319 ( .A1(n5893), .A2(n6168), .B1(n5117), .B2(n6454), .C1(n6167), 
        .C2(\intadd_2/SUM[4] ), .ZN(btb_cache_data_in[5]) );
  OAI222_X1 U7320 ( .A1(n5881), .A2(n6168), .B1(n5117), .B2(n6457), .C1(n3870), 
        .C2(\intadd_2/SUM[3] ), .ZN(btb_cache_data_in[4]) );
  OAI222_X1 U7321 ( .A1(n5864), .A2(n6168), .B1(n5117), .B2(n6460), .C1(n6167), 
        .C2(\intadd_2/SUM[2] ), .ZN(btb_cache_data_in[3]) );
  OAI222_X1 U7322 ( .A1(n5850), .A2(n6168), .B1(n5117), .B2(n6462), .C1(n3870), 
        .C2(\intadd_2/SUM[1] ), .ZN(btb_cache_data_in[2]) );
  OAI222_X1 U7323 ( .A1(n5836), .A2(n6168), .B1(n5117), .B2(n6464), .C1(n6167), 
        .C2(\intadd_2/SUM[0] ), .ZN(btb_cache_data_in[1]) );
  OAI222_X1 U7324 ( .A1(n6114), .A2(n6168), .B1(n5117), .B2(n6414), .C1(n3870), 
        .C2(\intadd_2/SUM[26] ), .ZN(btb_cache_data_in[27]) );
  OAI211_X1 U7325 ( .C1(alu_comp_sel[0]), .C2(n7086), .A(n7085), .B(
        alu_comp_sel[1]), .ZN(n7088) );
  NAND2_X1 U7326 ( .A1(\intadd_1/A[0] ), .A2(\intadd_1/B[0] ), .ZN(
        \intadd_1/n172 ) );
  NOR2_X1 U7327 ( .A1(\intadd_1/A[0] ), .A2(\intadd_1/B[0] ), .ZN(
        \intadd_1/n171 ) );
  NAND2_X1 U7328 ( .A1(n3897), .A2(\dp/b_mult_id_exe_int[2] ), .ZN(n6900) );
  NAND2_X1 U7329 ( .A1(n5211), .A2(\dp/b_mult_id_exe_int[2] ), .ZN(n6898) );
  NOR3_X1 U7330 ( .A1(\dp/b_mult_id_exe_int[2] ), .A2(n594), .A3(n595), .ZN(
        n5687) );
  NAND2_X1 U7331 ( .A1(n3900), .A2(\dp/b_mult_id_exe_int[2] ), .ZN(n5686) );
  NAND2_X1 U7332 ( .A1(n7256), .A2(n5262), .ZN(n5828) );
  XNOR2_X1 U7333 ( .A(rt_id[0]), .B(rd_exemem[0]), .ZN(n5366) );
  XNOR2_X1 U7334 ( .A(n4019), .B(n4083), .ZN(n5357) );
  AOI21_X1 U7335 ( .B1(n5122), .B2(\dp/b_adder_id_exe_int[4] ), .A(n7254), 
        .ZN(n5837) );
  NAND2_X1 U7336 ( .A1(n5120), .A2(n4345), .ZN(n5247) );
  NAND2_X1 U7337 ( .A1(n5120), .A2(n4346), .ZN(n5249) );
  NAND2_X1 U7338 ( .A1(\intadd_1/A[8] ), .A2(\intadd_1/B[8] ), .ZN(
        \intadd_1/n135 ) );
  XNOR2_X1 U7339 ( .A(n5828), .B(sub_add_exe), .ZN(\intadd_1/A[2] ) );
  AND2_X1 U7340 ( .A1(n5684), .A2(n3900), .ZN(n5153) );
  NOR2_X1 U7341 ( .A1(n5680), .A2(n5679), .ZN(n5684) );
  OAI21_X1 U7342 ( .B1(n5670), .B2(n4595), .A(n5233), .ZN(\ctrl_u/n559 ) );
  AOI21_X1 U7343 ( .B1(n5670), .B2(\ctrl_u/curr_mul_end_mem ), .A(n5229), .ZN(
        n5233) );
  AOI22_X1 U7344 ( .A1(n5670), .A2(\ctrl_u/curr_exe[6] ), .B1(n7340), .B2(
        \ctrl_u/curr_mem[6] ), .ZN(n5664) );
  AOI22_X1 U7345 ( .A1(n5670), .A2(\ctrl_u/curr_exe[4] ), .B1(n7340), .B2(
        \ctrl_u/curr_mem[4] ), .ZN(n5663) );
  AOI22_X1 U7346 ( .A1(n5670), .A2(\ctrl_u/curr_exe[2] ), .B1(n7340), .B2(
        \ctrl_u/curr_mem[2] ), .ZN(n5661) );
  AOI22_X1 U7347 ( .A1(n5670), .A2(\ctrl_u/curr_exe[3] ), .B1(
        \ctrl_u/curr_mem[3] ), .B2(n7340), .ZN(n5662) );
  OAI21_X1 U7348 ( .B1(n5654), .B2(n5659), .A(n5670), .ZN(\ctrl_u/exe_stall )
         );
  OR3_X1 U7349 ( .A1(n5658), .A2(wr_mem), .A3(n5341), .ZN(n5769) );
  NOR2_X1 U7350 ( .A1(n4038), .A2(\intadd_1/B[10] ), .ZN(\intadd_1/n122 ) );
  NAND2_X1 U7351 ( .A1(\intadd_1/A[11] ), .A2(\intadd_1/B[11] ), .ZN(
        \intadd_1/n115 ) );
  AOI22_X1 U7352 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[63] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[63] ), .ZN(n6325) );
  AOI22_X1 U7353 ( .A1(n3939), .A2(\dp/a_neg_mult_id_exe_int[24] ), .B1(n5185), 
        .B2(\dp/a_mult_id_exe_int[24] ), .ZN(n6045) );
  NAND2_X1 U7354 ( .A1(n5684), .A2(n5682), .ZN(n5683) );
  NAND2_X1 U7355 ( .A1(n5684), .A2(n3899), .ZN(n5712) );
  NOR2_X1 U7356 ( .A1(n5659), .A2(n5658), .ZN(n5669) );
  NAND2_X1 U7357 ( .A1(\intadd_1/A[7] ), .A2(\intadd_1/B[7] ), .ZN(
        \intadd_1/n138 ) );
  NOR2_X1 U7358 ( .A1(n5683), .A2(n4231), .ZN(n6322) );
  AOI22_X1 U7359 ( .A1(n6323), .A2(\dp/a_neg_mult_id_exe_int[1] ), .B1(n6322), 
        .B2(\dp/a_mult_id_exe_int[2] ), .ZN(n5718) );
  NAND2_X1 U7360 ( .A1(n5120), .A2(\dp/b_adder_id_exe_int[2] ), .ZN(n5323) );
  NAND2_X1 U7361 ( .A1(n5156), .A2(\dp/mul_feedback_exe_mem_int[1] ), .ZN(
        n5716) );
  XNOR2_X1 U7362 ( .A(\intadd_1/n89 ), .B(\intadd_1/n11 ), .ZN(
        \intadd_1/SUM[15] ) );
  AOI21_X1 U7363 ( .B1(\intadd_1/n89 ), .B2(\intadd_1/n85 ), .A(\intadd_1/n86 ), .ZN(\intadd_1/n84 ) );
  OAI21_X1 U7364 ( .B1(\intadd_1/n150 ), .B2(\intadd_1/n148 ), .A(
        \intadd_1/n149 ), .ZN(\intadd_1/n147 ) );
  OAI21_X1 U7365 ( .B1(\intadd_1/n145 ), .B2(\intadd_1/n149 ), .A(
        \intadd_1/n146 ), .ZN(\intadd_1/n144 ) );
  XNOR2_X1 U7366 ( .A(n5882), .B(sub_add_exe), .ZN(\intadd_1/A[6] ) );
  OAI21_X1 U7367 ( .B1(\intadd_1/n169 ), .B2(n3905), .A(\intadd_1/n168 ), .ZN(
        \intadd_1/n166 ) );
  NAND2_X1 U7368 ( .A1(\intadd_1/n198 ), .A2(\intadd_1/n168 ), .ZN(
        \intadd_1/n25 ) );
  NAND2_X1 U7369 ( .A1(\intadd_1/A[12] ), .A2(\intadd_1/B[12] ), .ZN(
        \intadd_1/n110 ) );
  NAND2_X1 U7370 ( .A1(n3903), .A2(\dp/b_adder_id_exe_int[3] ), .ZN(n5262) );
  INV_X1 U7371 ( .A(n5814), .ZN(n5815) );
  NAND2_X1 U7372 ( .A1(n6467), .A2(n6468), .ZN(n6466) );
  OAI211_X1 U7373 ( .C1(n3960), .C2(n4239), .A(n5717), .B(n5716), .ZN(n6467)
         );
  AOI21_X1 U7374 ( .B1(\intadd_1/n143 ), .B2(\intadd_1/n152 ), .A(
        \intadd_1/n144 ), .ZN(\intadd_1/n142 ) );
  NAND2_X1 U7375 ( .A1(n5120), .A2(n4347), .ZN(n5255) );
  AOI21_X1 U7376 ( .B1(n5122), .B2(n4343), .A(n5242), .ZN(n6036) );
  NAND2_X1 U7377 ( .A1(n5119), .A2(n4348), .ZN(n5258) );
  OAI21_X1 U7378 ( .B1(n5736), .B2(n5735), .A(n5897), .ZN(n5737) );
  AND2_X1 U7379 ( .A1(n5354), .A2(n5164), .ZN(n5356) );
  NAND2_X1 U7380 ( .A1(n5164), .A2(n5162), .ZN(n5348) );
  INV_X1 U7381 ( .A(n5732), .ZN(n5736) );
  OAI21_X1 U7382 ( .B1(\intadd_1/n122 ), .B2(\intadd_1/n128 ), .A(
        \intadd_1/n123 ), .ZN(\intadd_1/n121 ) );
  AOI21_X1 U7383 ( .B1(\intadd_1/n95 ), .B2(\intadd_1/n108 ), .A(
        \intadd_1/n96 ), .ZN(\intadd_1/n94 ) );
  OAI21_X1 U7384 ( .B1(\intadd_1/n103 ), .B2(\intadd_1/n97 ), .A(
        \intadd_1/n98 ), .ZN(\intadd_1/n96 ) );
  OAI21_X1 U7385 ( .B1(\intadd_1/n115 ), .B2(\intadd_1/n109 ), .A(
        \intadd_1/n110 ), .ZN(\intadd_1/n108 ) );
  NAND2_X1 U7386 ( .A1(\intadd_1/n85 ), .A2(\intadd_1/n88 ), .ZN(
        \intadd_1/n11 ) );
  OAI21_X1 U7387 ( .B1(\intadd_1/n82 ), .B2(\intadd_1/n88 ), .A(\intadd_1/n83 ), .ZN(\intadd_1/n81 ) );
  NOR2_X1 U7388 ( .A1(\intadd_1/A[15] ), .A2(\intadd_1/B[15] ), .ZN(
        \intadd_1/n87 ) );
  NAND2_X1 U7389 ( .A1(\intadd_1/A[15] ), .A2(\intadd_1/B[15] ), .ZN(
        \intadd_1/n88 ) );
  OAI21_X1 U7390 ( .B1(\intadd_1/n53 ), .B2(\intadd_1/n57 ), .A(\intadd_1/n54 ), .ZN(\intadd_1/n52 ) );
  NAND2_X1 U7391 ( .A1(\intadd_1/A[21] ), .A2(\intadd_1/B[21] ), .ZN(
        \intadd_1/n57 ) );
  AOI21_X1 U7392 ( .B1(\intadd_1/n51 ), .B2(\intadd_1/n60 ), .A(\intadd_1/n52 ), .ZN(\intadd_1/n50 ) );
  OAI21_X1 U7393 ( .B1(n4026), .B2(\intadd_1/n65 ), .A(\intadd_1/n62 ), .ZN(
        \intadd_1/n60 ) );
  NAND2_X1 U7394 ( .A1(\intadd_1/A[18] ), .A2(\intadd_1/B[18] ), .ZN(
        \intadd_1/n75 ) );
  OAI21_X1 U7395 ( .B1(\intadd_1/n74 ), .B2(\intadd_1/n78 ), .A(\intadd_1/n75 ), .ZN(\intadd_1/n73 ) );
  AOI21_X1 U7396 ( .B1(n5885), .B2(n5886), .A(n5898), .ZN(n5733) );
  XNOR2_X1 U7397 ( .A(n5898), .B(n5897), .ZN(n5899) );
  NAND2_X1 U7398 ( .A1(n5725), .A2(n5726), .ZN(n5166) );
  AOI21_X1 U7399 ( .B1(n5698), .B2(n5872), .A(n5697), .ZN(n5726) );
  NAND2_X1 U7400 ( .A1(\intadd_1/A[14] ), .A2(\intadd_1/B[14] ), .ZN(
        \intadd_1/n98 ) );
  OAI22_X1 U7401 ( .A1(n5132), .A2(n7129), .B1(n380), .B2(n4850), .ZN(n3020)
         );
  NAND2_X1 U7402 ( .A1(\intadd_1/B[1] ), .A2(\intadd_1/A[1] ), .ZN(
        \intadd_1/n168 ) );
  NAND2_X1 U7403 ( .A1(n5739), .A2(n5738), .ZN(n5919) );
  OAI21_X1 U7404 ( .B1(sub_add_exe), .B2(n7071), .A(n5328), .ZN(\intadd_1/CI )
         );
  NAND2_X1 U7405 ( .A1(n7064), .A2(n7071), .ZN(n5328) );
  NAND2_X1 U7406 ( .A1(n5900), .A2(n5898), .ZN(n5167) );
  NAND2_X1 U7407 ( .A1(n5167), .A2(n5737), .ZN(n5911) );
  XNOR2_X1 U7408 ( .A(n5900), .B(n5899), .ZN(n5901) );
  OAI211_X1 U7409 ( .C1(n3920), .C2(alu_comp_sel[0]), .A(n7092), .B(n4139), 
        .ZN(n7093) );
  NAND2_X1 U7410 ( .A1(n5731), .A2(n5732), .ZN(n5900) );
  NAND2_X1 U7411 ( .A1(n5730), .A2(n5886), .ZN(n5731) );
  OR2_X1 U7412 ( .A1(n5348), .A2(n5148), .ZN(n5351) );
  NAND2_X1 U7413 ( .A1(\dp/exs/alu_unit/mult/ax2_shiftn[4] ), .A2(n6298), .ZN(
        n5704) );
  OAI22_X1 U7414 ( .A1(n5584), .A2(n5569), .B1(n5182), .B2(n4396), .ZN(
        \ctrl_u/n554 ) );
  NAND2_X1 U7415 ( .A1(n4038), .A2(\intadd_1/B[10] ), .ZN(\intadd_1/n123 ) );
  OAI21_X1 U7416 ( .B1(n5166), .B2(n5734), .A(n5733), .ZN(n5735) );
  NAND2_X1 U7417 ( .A1(n5166), .A2(n5729), .ZN(n5730) );
  XNOR2_X1 U7418 ( .A(n5888), .B(n5887), .ZN(n5889) );
  NAND2_X1 U7419 ( .A1(n5888), .A2(n5885), .ZN(n5732) );
  AOI21_X1 U7420 ( .B1(\intadd_1/n89 ), .B2(\intadd_1/n47 ), .A(\intadd_1/n48 ), .ZN(\intadd_1/n46 ) );
  OAI211_X1 U7421 ( .C1(n5840), .C2(n5841), .A(n5720), .B(n5842), .ZN(n5723)
         );
  AOI21_X1 U7422 ( .B1(\dp/exs/alu_unit/mult/neg_ax2_shiftn[4] ), .B2(n6326), 
        .A(n5703), .ZN(n5705) );
  OAI21_X1 U7423 ( .B1(n3882), .B2(n5165), .A(n5353), .ZN(\ctrl_u/n503 ) );
  AND2_X1 U7424 ( .A1(n7274), .A2(n5165), .ZN(n5352) );
  INV_X1 U7425 ( .A(n5701), .ZN(n5698) );
  NAND2_X1 U7426 ( .A1(n5701), .A2(n5700), .ZN(n5724) );
  NAND2_X1 U7427 ( .A1(\dp/exs/alu_unit/mult/ax2_shiftn[6] ), .A2(n6298), .ZN(
        n5690) );
  OAI21_X1 U7428 ( .B1(n5493), .B2(n5492), .A(n5510), .ZN(n5539) );
  INV_X1 U7429 ( .A(n5510), .ZN(n5584) );
  OAI22_X1 U7430 ( .A1(n6412), .A2(n7440), .B1(n4109), .B2(n3938), .ZN(n2623)
         );
  INV_X1 U7431 ( .A(n6412), .ZN(n6413) );
  OAI211_X1 U7432 ( .C1(n6119), .C2(n6141), .A(n6118), .B(n6117), .ZN(n6120)
         );
  INV_X1 U7433 ( .A(n6119), .ZN(n6116) );
  NAND2_X1 U7434 ( .A1(n6119), .A2(n6141), .ZN(n6122) );
  XNOR2_X1 U7435 ( .A(n5957), .B(n5759), .ZN(n5766) );
  AOI21_X1 U7436 ( .B1(n5870), .B2(n5869), .A(n5868), .ZN(n5871) );
  INV_X1 U7437 ( .A(n5868), .ZN(n5694) );
  NAND2_X1 U7438 ( .A1(\dp/exs/alu_unit/mult/ax2_shiftn[5] ), .A2(n5187), .ZN(
        n5707) );
  XNOR2_X1 U7439 ( .A(n6055), .B(n6046), .ZN(n6053) );
  AOI21_X1 U7440 ( .B1(\dp/exs/alu_unit/mult/neg_ax2_shiftn[6] ), .B2(n6326), 
        .A(n5689), .ZN(n5691) );
  OAI22_X1 U7441 ( .A1(n3927), .A2(n5517), .B1(n5182), .B2(n4600), .ZN(
        \ctrl_u/n526 ) );
  NOR2_X1 U7442 ( .A1(n5653), .A2(n5526), .ZN(n5527) );
  NOR2_X1 U7443 ( .A1(n3927), .A2(n5521), .ZN(n5528) );
  OAI211_X1 U7444 ( .C1(\intadd_1/SUM[14] ), .C2(n7066), .A(n5949), .B(n5948), 
        .ZN(n5950) );
  OAI21_X1 U7445 ( .B1(\intadd_1/n139 ), .B2(\intadd_1/n137 ), .A(
        \intadd_1/n138 ), .ZN(\intadd_1/n136 ) );
  XOR2_X1 U7446 ( .A(\intadd_1/n139 ), .B(\intadd_1/n19 ), .Z(
        \intadd_1/SUM[7] ) );
  NOR2_X1 U7447 ( .A1(\intadd_1/n164 ), .A2(\intadd_1/n167 ), .ZN(
        \intadd_1/n162 ) );
  OAI21_X1 U7448 ( .B1(\intadd_1/n168 ), .B2(\intadd_1/n164 ), .A(
        \intadd_1/n165 ), .ZN(\intadd_1/n163 ) );
  NAND2_X1 U7449 ( .A1(n7274), .A2(n5155), .ZN(n5346) );
  NAND2_X1 U7450 ( .A1(n3911), .A2(n5719), .ZN(n5720) );
  OAI21_X1 U7451 ( .B1(n5858), .B2(n3911), .A(n5857), .ZN(n5870) );
  OAI22_X1 U7452 ( .A1(n6621), .A2(n7062), .B1(n4194), .B2(n3938), .ZN(n2799)
         );
  XNOR2_X1 U7453 ( .A(n5969), .B(n5960), .ZN(n5967) );
  NAND2_X1 U7454 ( .A1(\dp/exs/alu_unit/mult/neg_ax2_shiftn[5] ), .A2(n5154), 
        .ZN(n5693) );
  NAND2_X1 U7455 ( .A1(\dp/exs/alu_unit/mult/neg_ax2_shiftn[5] ), .A2(n5188), 
        .ZN(n5706) );
  XNOR2_X1 U7456 ( .A(n3917), .B(n6081), .ZN(n6086) );
  NAND2_X1 U7457 ( .A1(n5699), .A2(n5872), .ZN(n5700) );
  NAND2_X1 U7458 ( .A1(n5699), .A2(n5694), .ZN(n5701) );
  NAND2_X1 U7459 ( .A1(n5655), .A2(n5418), .ZN(n5674) );
  OAI22_X1 U7460 ( .A1(n4040), .A2(wp_data[26]), .B1(
        \dp/mul_feedback_exe_mem_int[26] ), .B2(n3922), .ZN(n5240) );
  OAI22_X1 U7461 ( .A1(n3913), .A2(wp_data[24]), .B1(
        \dp/mul_feedback_exe_mem_int[24] ), .B2(n3922), .ZN(n5241) );
  OAI22_X1 U7462 ( .A1(n4040), .A2(wp_data[14]), .B1(
        \dp/mul_feedback_exe_mem_int[14] ), .B2(n3922), .ZN(n5250) );
  OAI21_X1 U7463 ( .B1(n3922), .B2(n4071), .A(n5261), .ZN(n7254) );
  OAI22_X1 U7464 ( .A1(n3913), .A2(wp_data[12]), .B1(
        \dp/mul_feedback_exe_mem_int[12] ), .B2(n3922), .ZN(n5252) );
  AOI22_X1 U7465 ( .A1(n5136), .A2(n4074), .B1(n5310), .B2(n4024), .ZN(n5254)
         );
  AOI22_X1 U7466 ( .A1(n5136), .A2(n4063), .B1(n5314), .B2(n4024), .ZN(n5257)
         );
  OAI22_X1 U7467 ( .A1(n4040), .A2(wp_data[22]), .B1(
        \dp/mul_feedback_exe_mem_int[22] ), .B2(n3922), .ZN(n5243) );
  AOI22_X1 U7468 ( .A1(n5136), .A2(n4081), .B1(n5301), .B2(n4024), .ZN(n5248)
         );
  OAI22_X1 U7469 ( .A1(n3913), .A2(wp_data[23]), .B1(
        \dp/mul_feedback_exe_mem_int[23] ), .B2(n3922), .ZN(n5242) );
  OAI22_X1 U7470 ( .A1(n5273), .A2(wp_data[6]), .B1(
        \dp/mul_feedback_exe_mem_int[6] ), .B2(n3922), .ZN(n5259) );
  OAI22_X1 U7471 ( .A1(n5273), .A2(wp_data[18]), .B1(
        \dp/mul_feedback_exe_mem_int[18] ), .B2(n3922), .ZN(n5245) );
  AOI22_X1 U7472 ( .A1(n5136), .A2(n4073), .B1(n5306), .B2(n3906), .ZN(n5253)
         );
  AOI22_X1 U7473 ( .A1(n5136), .A2(n4095), .B1(n5295), .B2(n4024), .ZN(n5246)
         );
  AOI22_X1 U7474 ( .A1(n5136), .A2(\dp/mul_feedback_exe_mem_int[2] ), .B1(
        n4024), .B2(wp_data[2]), .ZN(n7257) );
  AOI22_X1 U7475 ( .A1(n5136), .A2(n4082), .B1(n5312), .B2(n4024), .ZN(n5256)
         );
  OAI22_X1 U7476 ( .A1(n4040), .A2(wp_data[19]), .B1(
        \dp/mul_feedback_exe_mem_int[19] ), .B2(n3922), .ZN(n5244) );
  OAI22_X1 U7477 ( .A1(n3913), .A2(wp_data[13]), .B1(n3922), .B2(
        \dp/mul_feedback_exe_mem_int[13] ), .ZN(n5251) );
  AOI22_X1 U7478 ( .A1(n4024), .A2(wp_data[0]), .B1(n5136), .B2(
        \dp/mul_feedback_exe_mem_int[0] ), .ZN(n7259) );
  OAI22_X1 U7479 ( .A1(n4040), .A2(wp_data[5]), .B1(
        \dp/mul_feedback_exe_mem_int[5] ), .B2(n3922), .ZN(n5260) );
  OAI22_X1 U7480 ( .A1(n5273), .A2(n5324), .B1(n3922), .B2(n4072), .ZN(n7258)
         );
  AOI22_X1 U7481 ( .A1(n5136), .A2(\dp/mul_feedback_exe_mem_int[3] ), .B1(
        n5140), .B2(wp_data[3]), .ZN(n7256) );
  XNOR2_X1 U7482 ( .A(n5931), .B(n5930), .ZN(n5937) );
  XNOR2_X1 U7483 ( .A(n6003), .B(n5994), .ZN(n6001) );
  XNOR2_X1 U7484 ( .A(n5945), .B(n5944), .ZN(n5951) );
  XNOR2_X1 U7485 ( .A(n4023), .B(n6104), .ZN(n6111) );
  OAI21_X1 U7486 ( .B1(n5158), .B2(n3882), .A(n5345), .ZN(\ctrl_u/n558 ) );
  OAI21_X1 U7487 ( .B1(n5545), .B2(n5544), .A(n5641), .ZN(n5546) );
  AOI22_X1 U7488 ( .A1(n5641), .A2(n5533), .B1(n3941), .B2(
        \ctrl_u/curr_id[28] ), .ZN(n5535) );
  OAI21_X1 U7489 ( .B1(n5134), .B2(n7186), .A(n5626), .ZN(n5429) );
  NAND2_X1 U7490 ( .A1(n5655), .A2(\ctrl_u/curr_id[29] ), .ZN(n5410) );
  AOI22_X1 U7491 ( .A1(n5407), .A2(\ctrl_u/curr_exe[18] ), .B1(n5655), .B2(
        \ctrl_u/curr_id[18] ), .ZN(n5400) );
  AOI22_X1 U7492 ( .A1(n5407), .A2(\ctrl_u/curr_exe[6] ), .B1(n5655), .B2(
        \ctrl_u/curr_id[6] ), .ZN(n5396) );
  AOI22_X1 U7493 ( .A1(n5407), .A2(\ctrl_u/curr_exe[4] ), .B1(n5655), .B2(
        \ctrl_u/curr_id[4] ), .ZN(n5394) );
  AOI22_X1 U7494 ( .A1(n5407), .A2(\ctrl_u/curr_exe[3] ), .B1(n5655), .B2(
        \ctrl_u/curr_id[3] ), .ZN(n5392) );
  AOI22_X1 U7495 ( .A1(n5407), .A2(\ctrl_u/curr_exe[2] ), .B1(n5655), .B2(
        \ctrl_u/curr_id[2] ), .ZN(n5390) );
  AOI22_X1 U7496 ( .A1(n5407), .A2(cond_sel_exe[2]), .B1(n5655), .B2(
        \ctrl_u/curr_id[26] ), .ZN(n5408) );
  AOI22_X1 U7497 ( .A1(n5407), .A2(alu_comp_sel[1]), .B1(n5655), .B2(
        \ctrl_u/curr_id[22] ), .ZN(n5402) );
  AND2_X1 U7498 ( .A1(n5655), .A2(n5618), .ZN(n5672) );
  NAND2_X1 U7499 ( .A1(n5160), .A2(\ctrl_u/n94 ), .ZN(n5168) );
  OAI22_X1 U7500 ( .A1(n6593), .A2(n7062), .B1(n4191), .B2(n3938), .ZN(n2803)
         );
  OAI22_X1 U7501 ( .A1(n6593), .A2(n5196), .B1(n4487), .B2(n5199), .ZN(n2835)
         );
  XNOR2_X1 U7502 ( .A(n3918), .B(n5910), .ZN(n5912) );
  XNOR2_X1 U7503 ( .A(n5874), .B(n5152), .ZN(n5875) );
  NAND2_X1 U7504 ( .A1(n5911), .A2(n5909), .ZN(n5738) );
  OAI21_X1 U7505 ( .B1(n5911), .B2(n5909), .A(n5908), .ZN(n5739) );
  NOR2_X1 U7506 ( .A1(n5874), .A2(n5152), .ZN(n5697) );
  NAND2_X1 U7507 ( .A1(n5874), .A2(n5152), .ZN(n5699) );
  AOI21_X1 U7508 ( .B1(n6714), .B2(n6695), .A(n6704), .ZN(n6697) );
  AOI21_X1 U7509 ( .B1(n3871), .B2(n6661), .A(n6665), .ZN(n6648) );
  AOI21_X1 U7510 ( .B1(n5124), .B2(n6713), .A(n6712), .ZN(n6718) );
  AOI21_X1 U7511 ( .B1(n3871), .B2(n6612), .A(n6614), .ZN(n6610) );
  AOI21_X1 U7512 ( .B1(n6714), .B2(n6486), .A(n6490), .ZN(n6484) );
  AOI21_X1 U7513 ( .B1(n5124), .B2(n6586), .A(n6588), .ZN(n6584) );
  AOI21_X1 U7514 ( .B1(n6714), .B2(n6622), .A(n6625), .ZN(n6595) );
  AOI21_X1 U7515 ( .B1(n5124), .B2(n6560), .A(n6563), .ZN(n6530) );
  AOI21_X1 U7516 ( .B1(n3871), .B2(n6480), .A(n6479), .ZN(n6481) );
  XNOR2_X1 U7517 ( .A(n6075), .B(n6064), .ZN(n6071) );
  XNOR2_X1 U7518 ( .A(n5988), .B(n5977), .ZN(n5984) );
  XNOR2_X1 U7519 ( .A(n6022), .B(n6011), .ZN(n6018) );
  XNOR2_X1 U7520 ( .A(n5855), .B(n5854), .ZN(n5845) );
  OAI21_X1 U7521 ( .B1(n5856), .B2(n5855), .A(n5854), .ZN(n5857) );
  NAND4_X1 U7522 ( .A1(n5724), .A2(n5723), .A3(n5722), .A4(n5721), .ZN(n5725)
         );
  NAND2_X1 U7523 ( .A1(n5855), .A2(n5854), .ZN(n5722) );
  INV_X1 U7524 ( .A(n5130), .ZN(n5180) );
  INV_X1 U7525 ( .A(\intadd_1/n102 ), .ZN(\intadd_1/n186 ) );
  INV_X1 U7526 ( .A(\intadd_1/n103 ), .ZN(\intadd_1/n101 ) );
  INV_X1 U7527 ( .A(\intadd_1/n114 ), .ZN(\intadd_1/n188 ) );
  INV_X1 U7528 ( .A(\intadd_1/n115 ), .ZN(\intadd_1/n113 ) );
  INV_X1 U7529 ( .A(\intadd_1/n127 ), .ZN(\intadd_1/n190 ) );
  INV_X1 U7530 ( .A(\intadd_1/n132 ), .ZN(\intadd_1/n130 ) );
  INV_X1 U7531 ( .A(\intadd_1/n158 ), .ZN(\intadd_1/n196 ) );
  INV_X1 U7532 ( .A(\intadd_1/n161 ), .ZN(\intadd_1/n160 ) );
  INV_X1 U7533 ( .A(n4029), .ZN(\intadd_1/n169 ) );
  INV_X1 U7534 ( .A(\intadd_1/CI ), .ZN(\intadd_1/n173 ) );
  INV_X1 U7535 ( .A(\intadd_1/n53 ), .ZN(\intadd_1/n177 ) );
  INV_X1 U7536 ( .A(n4026), .ZN(\intadd_1/n179 ) );
  INV_X1 U7537 ( .A(n3861), .ZN(\intadd_1/n181 ) );
  INV_X1 U7538 ( .A(\intadd_1/n77 ), .ZN(\intadd_1/n182 ) );
  INV_X1 U7539 ( .A(\intadd_1/n82 ), .ZN(\intadd_1/n183 ) );
  INV_X1 U7540 ( .A(\intadd_1/n87 ), .ZN(\intadd_1/n85 ) );
  INV_X1 U7541 ( .A(n3916), .ZN(\intadd_1/n185 ) );
  INV_X1 U7542 ( .A(\intadd_1/n134 ), .ZN(\intadd_1/n191 ) );
  INV_X1 U7543 ( .A(\intadd_1/n137 ), .ZN(\intadd_1/n192 ) );
  INV_X1 U7544 ( .A(\intadd_1/n145 ), .ZN(\intadd_1/n193 ) );
  INV_X1 U7545 ( .A(\intadd_1/n167 ), .ZN(\intadd_1/n198 ) );
  INV_X1 U7546 ( .A(\intadd_1/n171 ), .ZN(\intadd_1/n199 ) );
  INV_X1 U7547 ( .A(\intadd_1/n45 ), .ZN(\intadd_1/n43 ) );
  INV_X1 U7548 ( .A(\intadd_1/n88 ), .ZN(\intadd_1/n86 ) );
  NAND3_X1 U7549 ( .A1(n6162), .A2(n6159), .A3(op_sign_exe), .ZN(n5335) );
  MUX2_X1 U7550 ( .A(n5354), .B(n5349), .S(n5164), .Z(\ctrl_u/n502 ) );
  NAND3_X1 U7551 ( .A1(n5621), .A2(n5352), .A3(n5351), .ZN(n5353) );
  MUX2_X1 U7552 ( .A(n5356), .B(n5355), .S(n5162), .Z(\ctrl_u/n501 ) );
  NAND3_X1 U7553 ( .A1(n5375), .A2(n5374), .A3(n5373), .ZN(n5384) );
  NAND3_X1 U7554 ( .A1(n5379), .A2(n5378), .A3(n5377), .ZN(n5383) );
  MUX2_X1 U7555 ( .A(n5424), .B(n4358), .S(n5626), .Z(n5426) );
  NAND3_X1 U7556 ( .A1(n5499), .A2(n5595), .A3(n5500), .ZN(n5577) );
  NAND3_X1 U7557 ( .A1(instr_if[28]), .A2(instr_if[29]), .A3(n5590), .ZN(n5522) );
  NAND3_X1 U7558 ( .A1(n5450), .A2(n5639), .A3(n5441), .ZN(n5442) );
  MUX2_X1 U7559 ( .A(n5442), .B(\ctrl_u/curr_id[22] ), .S(n5626), .Z(n5443) );
  MUX2_X1 U7560 ( .A(n5453), .B(n4491), .S(n5626), .Z(n5454) );
  NAND3_X1 U7561 ( .A1(n5499), .A2(instr_if[4]), .A3(n5455), .ZN(n5456) );
  MUX2_X1 U7562 ( .A(n5472), .B(\ctrl_u/n61 ), .S(n5626), .Z(n5473) );
  NAND3_X1 U7563 ( .A1(n5475), .A2(n5474), .A3(n5522), .ZN(n5476) );
  MUX2_X1 U7564 ( .A(n5478), .B(\ctrl_u/n59 ), .S(n5626), .Z(n5479) );
  NAND3_X1 U7565 ( .A1(n5641), .A2(n5579), .A3(n7280), .ZN(n5484) );
  NAND3_X1 U7566 ( .A1(n5641), .A2(instr_if[1]), .A3(n5579), .ZN(n5486) );
  NAND3_X1 U7567 ( .A1(instr_if[30]), .A2(n5591), .A3(n7276), .ZN(n5512) );
  NAND3_X1 U7568 ( .A1(instr_if[3]), .A2(n5541), .A3(n5498), .ZN(n5624) );
  NAND3_X1 U7569 ( .A1(n5560), .A2(n5590), .A3(n5644), .ZN(n5503) );
  NAND3_X1 U7570 ( .A1(n5535), .A2(n5536), .A3(n5571), .ZN(\ctrl_u/n531 ) );
  NAND3_X1 U7571 ( .A1(n5641), .A2(n5602), .A3(n5601), .ZN(n5603) );
  MUX2_X1 U7572 ( .A(n5612), .B(\ctrl_u/n70 ), .S(n5626), .Z(n5613) );
  MUX2_X1 U7573 ( .A(n5614), .B(n4484), .S(n5626), .Z(n5615) );
  NAND3_X1 U7574 ( .A1(n5641), .A2(n5640), .A3(n5639), .ZN(n5642) );
  NAND3_X1 U7575 ( .A1(n5672), .A2(n5671), .A3(n5670), .ZN(n5673) );
  NAND3_X1 U7576 ( .A1(n5720), .A2(n5840), .A3(n5841), .ZN(n5721) );
  FA_X1 U7577 ( .A(n5917), .B(n5918), .CI(n5919), .CO(n5923) );
  MUX2_X1 U7578 ( .A(n7069), .B(n7080), .S(n5760), .Z(n5762) );
  MUX2_X1 U7579 ( .A(n5762), .B(n5761), .S(\intadd_1/B[16] ), .Z(n5763) );
  MUX2_X1 U7580 ( .A(n5813), .B(n5812), .S(\intadd_1/A[1] ), .Z(n5819) );
  MUX2_X1 U7581 ( .A(n7080), .B(n7069), .S(n5828), .Z(n5830) );
  MUX2_X1 U7582 ( .A(n5830), .B(n5829), .S(\intadd_1/B[2] ), .Z(n5834) );
  MUX2_X1 U7583 ( .A(n7069), .B(n6157), .S(\intadd_1/B[3] ), .Z(n5839) );
  MUX2_X1 U7584 ( .A(n5839), .B(n5838), .S(n5837), .Z(n5848) );
  MUX2_X1 U7585 ( .A(n7080), .B(n7069), .S(n5851), .Z(n5853) );
  MUX2_X1 U7586 ( .A(n5853), .B(n5852), .S(\intadd_1/B[4] ), .Z(n5862) );
  XOR2_X1 U7587 ( .A(n5872), .B(n5868), .Z(n5859) );
  MUX2_X1 U7588 ( .A(n7080), .B(n7069), .S(n5865), .Z(n5867) );
  MUX2_X1 U7589 ( .A(n5867), .B(n5866), .S(\intadd_1/B[5] ), .Z(n5879) );
  MUX2_X1 U7590 ( .A(n7080), .B(n7069), .S(n4042), .Z(n5884) );
  MUX2_X1 U7591 ( .A(n5884), .B(n5883), .S(\intadd_1/B[6] ), .Z(n5891) );
  MUX2_X1 U7592 ( .A(n7069), .B(n7080), .S(n5894), .Z(n5896) );
  MUX2_X1 U7593 ( .A(n5896), .B(n5895), .S(\intadd_1/B[7] ), .Z(n5903) );
  MUX2_X1 U7594 ( .A(n7069), .B(n7080), .S(n4672), .Z(n5907) );
  MUX2_X1 U7595 ( .A(n5907), .B(n5906), .S(\intadd_1/B[8] ), .Z(n5914) );
  XOR2_X1 U7596 ( .A(n5929), .B(n5928), .Z(n5930) );
  MUX2_X1 U7597 ( .A(n5933), .B(n5932), .S(\intadd_1/B[12] ), .Z(n5934) );
  MUX2_X1 U7598 ( .A(n5947), .B(n5946), .S(\intadd_1/B[14] ), .Z(n5949) );
  XOR2_X1 U7599 ( .A(n5971), .B(n5970), .Z(n5960) );
  MUX2_X1 U7600 ( .A(n7080), .B(n7069), .S(n5961), .Z(n5963) );
  MUX2_X1 U7601 ( .A(n5963), .B(n5962), .S(\intadd_1/B[17] ), .Z(n5964) );
  XOR2_X1 U7602 ( .A(n5986), .B(n5987), .Z(n5977) );
  MUX2_X1 U7603 ( .A(n7080), .B(n7069), .S(n5978), .Z(n5980) );
  MUX2_X1 U7604 ( .A(n5980), .B(n5979), .S(\intadd_1/B[18] ), .Z(n5981) );
  XOR2_X1 U7605 ( .A(n6005), .B(n6004), .Z(n5994) );
  MUX2_X1 U7606 ( .A(n7080), .B(n7069), .S(n5995), .Z(n5997) );
  MUX2_X1 U7607 ( .A(n5997), .B(n5996), .S(\intadd_1/B[19] ), .Z(n5998) );
  XOR2_X1 U7608 ( .A(n6020), .B(n6021), .Z(n6011) );
  MUX2_X1 U7609 ( .A(n7080), .B(n7069), .S(n6012), .Z(n6014) );
  MUX2_X1 U7610 ( .A(n6014), .B(n6013), .S(\intadd_1/B[20] ), .Z(n6015) );
  MUX2_X1 U7611 ( .A(n7080), .B(n7069), .S(n6036), .Z(n6037) );
  MUX2_X1 U7612 ( .A(n7080), .B(n7069), .S(n6047), .Z(n6049) );
  MUX2_X1 U7613 ( .A(n6049), .B(n6048), .S(\intadd_1/B[23] ), .Z(n6050) );
  FA_X1 U7614 ( .A(n6057), .B(n6056), .CI(n6055), .CO(n6075) );
  MUX2_X1 U7615 ( .A(n7069), .B(n7080), .S(n6065), .Z(n6067) );
  MUX2_X1 U7616 ( .A(n6067), .B(n6066), .S(\intadd_1/B[24] ), .Z(n6068) );
  MUX2_X1 U7617 ( .A(n7069), .B(n7080), .S(n6105), .Z(n6107) );
  MUX2_X1 U7618 ( .A(n6107), .B(n6106), .S(\intadd_1/B[27] ), .Z(n6109) );
  MUX2_X1 U7619 ( .A(n7069), .B(n7080), .S(n6124), .Z(n6126) );
  MUX2_X1 U7620 ( .A(n6126), .B(n6125), .S(\intadd_1/B[29] ), .Z(n6128) );
  XOR2_X1 U7621 ( .A(n6306), .B(n6307), .Z(n6156) );
  NAND3_X1 U7622 ( .A1(n6169), .A2(btb_cache_data_out_rw[31]), .A3(taken), 
        .ZN(n6170) );
  XOR2_X1 U7623 ( .A(n6330), .B(n6329), .Z(n6331) );
  XOR2_X1 U7624 ( .A(n6516), .B(n6515), .Z(n6517) );
  XOR2_X1 U7625 ( .A(n6545), .B(n6544), .Z(n6546) );
  XOR2_X1 U7626 ( .A(n6565), .B(n6564), .Z(n6566) );
  XOR2_X1 U7627 ( .A(n6627), .B(n6626), .Z(n6628) );
  XOR2_X1 U7628 ( .A(n6667), .B(n6666), .Z(n6668) );
  NAND3_X1 U7629 ( .A1(sign_ext_sel_id), .A2(is_signed_id), .A3(
        \dp/imm_id_int[15] ), .ZN(n7146) );
  NAND3_X1 U7630 ( .A1(n6963), .A2(n6925), .A3(n6924), .ZN(n2690) );
  NAND3_X1 U7631 ( .A1(n6963), .A2(n6927), .A3(n6926), .ZN(n2688) );
  NAND3_X1 U7632 ( .A1(n6963), .A2(n6960), .A3(n6959), .ZN(n2691) );
  NAND3_X1 U7633 ( .A1(n6963), .A2(n6962), .A3(n6961), .ZN(n2689) );
  MUX2_X1 U7634 ( .A(\dp/a_mult_id_exe_int[0] ), .B(
        \dp/mul_feedback_exe_mem_int[0] ), .S(n5186), .Z(n7072) );
  MUX2_X1 U7635 ( .A(n7072), .B(\dp/a_neg_mult_id_exe_int[0] ), .S(n3939), .Z(
        n7073) );
  NAND3_X1 U7636 ( .A1(n3932), .A2(en_rd_id), .A3(n4396), .ZN(n7165) );
  NAND3_X1 U7637 ( .A1(n3932), .A2(j_instr_id), .A3(en_rd_id), .ZN(n7168) );
  NOR2_X1 U7638 ( .A1(\ctrl_u/if_stall ), .A2(n4547), .ZN(\ctrl_u/n9 ) );
  NOR2_X1 U7639 ( .A1(\ctrl_u/if_stall ), .A2(\ctrl_u/n62 ), .ZN(\ctrl_u/n11 )
         );
  NOR2_X1 U7640 ( .A1(\ctrl_u/if_stall ), .A2(\ctrl_u/n64 ), .ZN(\ctrl_u/n13 )
         );
  NOR2_X1 U7641 ( .A1(\ctrl_u/if_stall ), .A2(\ctrl_u/n63 ), .ZN(\ctrl_u/n15 )
         );
  NOR2_X1 U7642 ( .A1(\ctrl_u/if_stall ), .A2(\ctrl_u/n65 ), .ZN(\ctrl_u/n21 )
         );
  NOR2_X1 U7643 ( .A1(\ctrl_u/if_stall ), .A2(\ctrl_u/n66 ), .ZN(\ctrl_u/n23 )
         );
  NOR2_X1 U7644 ( .A1(\ctrl_u/if_stall ), .A2(\ctrl_u/n67 ), .ZN(\ctrl_u/n25 )
         );
  NOR2_X1 U7645 ( .A1(\ctrl_u/if_stall ), .A2(\ctrl_u/n68 ), .ZN(\ctrl_u/n27 )
         );
  NOR2_X1 U7646 ( .A1(instr_if[3]), .A2(instr_if[2]), .ZN(n7288) );
  AOI221_X1 U7647 ( .B1(instr_if[2]), .B2(n7279), .C1(n7287), .C2(n7279), .A(
        n7290), .ZN(n7289) );
  OAI211_X1 U7648 ( .C1(n7291), .C2(n7281), .A(n7286), .B(n7285), .ZN(n7290)
         );
  AOI211_X1 U7649 ( .C1(n7283), .C2(n7287), .A(n7292), .B(n7282), .ZN(n7286)
         );
  OAI211_X1 U7650 ( .C1(instr_if[1]), .C2(n7291), .A(n7293), .B(n7294), .ZN(
        n7282) );
  NAND3_X1 U7651 ( .A1(instr_if[5]), .A2(instr_if[4]), .A3(n7279), .ZN(n7294)
         );
  AOI221_X1 U7652 ( .B1(n7264), .B2(n7277), .C1(n7284), .C2(instr_if[5]), .A(
        n7278), .ZN(n7292) );
  NOR2_X1 U7653 ( .A1(instr_if[2]), .A2(n7280), .ZN(n7283) );
  AOI221_X1 U7654 ( .B1(n7277), .B2(n7278), .C1(n7281), .C2(n7278), .A(
        instr_if[2]), .ZN(n7295) );
  NAND2_X1 U7655 ( .A1(n7277), .A2(instr_if[2]), .ZN(n7291) );
  NOR2_X1 U7656 ( .A1(n7276), .A2(n7275), .ZN(n7296) );
  NOR2_X1 U7657 ( .A1(instr_if[5]), .A2(instr_if[4]), .ZN(n7287) );
  NOR2_X1 U7658 ( .A1(instr_if[9]), .A2(n7297), .ZN(n7293) );
  OR4_X1 U7659 ( .A1(instr_if[10]), .A2(instr_if[6]), .A3(instr_if[7]), .A4(
        instr_if[8]), .ZN(n7297) );
  INV_X1 U7660 ( .A(\ctrl_u/exe_stall ), .ZN(n7298) );
  NOR2_X1 U7661 ( .A1(\ctrl_u/next_mem[2] ), .A2(n5229), .ZN(\ctrl_u/n478 ) );
  NOR2_X1 U7662 ( .A1(\ctrl_u/next_mem[3] ), .A2(n5229), .ZN(\ctrl_u/n477 ) );
  NOR2_X1 U7663 ( .A1(\ctrl_u/next_mem[4] ), .A2(n5229), .ZN(\ctrl_u/n476 ) );
  NOR2_X1 U7664 ( .A1(\ctrl_u/next_mem[6] ), .A2(n5229), .ZN(\ctrl_u/n474 ) );
  NAND2_X1 U7665 ( .A1(rst_mem_wb_regs), .A2(\ctrl_u/next_mem[7] ), .ZN(
        \ctrl_u/n473 ) );
  NAND2_X1 U7666 ( .A1(rst_mem_wb_regs), .A2(\ctrl_u/next_mem[8] ), .ZN(
        \ctrl_u/n472 ) );
  NAND2_X1 U7667 ( .A1(rst_mem_wb_regs), .A2(\ctrl_u/next_mem[10] ), .ZN(
        \ctrl_u/n470 ) );
  NOR2_X1 U7668 ( .A1(n5158), .A2(n4025), .ZN(\ctrl_u/N1805 ) );
  OAI22_X1 U7670 ( .A1(n4138), .A2(rd_idexe[1]), .B1(n4365), .B2(rd_idexe[2]), 
        .ZN(n7299) );
  AOI221_X1 U7671 ( .B1(n4138), .B2(rd_idexe[1]), .C1(rd_idexe[2]), .C2(n4365), 
        .A(n7299), .ZN(n7303) );
  OAI22_X1 U7672 ( .A1(n4212), .A2(rd_idexe[3]), .B1(n4240), .B2(rt_id[0]), 
        .ZN(n7300) );
  AOI221_X1 U7673 ( .B1(n4212), .B2(rd_idexe[3]), .C1(rt_id[0]), .C2(n4240), 
        .A(n7300), .ZN(n7302) );
  XOR2_X1 U7674 ( .A(n4359), .B(rd_idexe[4]), .Z(n7301) );
  NAND4_X1 U7675 ( .A1(\ctrl_u/curr_exe[15] ), .A2(n7303), .A3(n7302), .A4(
        n7301), .ZN(n7311) );
  OAI22_X1 U7676 ( .A1(rd_idexe[3]), .A2(n4366), .B1(n4370), .B2(rd_idexe[2]), 
        .ZN(n7304) );
  AOI221_X1 U7677 ( .B1(n4366), .B2(rd_idexe[3]), .C1(n4370), .C2(rd_idexe[2]), 
        .A(n7304), .ZN(n7308) );
  OAI22_X1 U7678 ( .A1(rd_idexe[0]), .A2(n4083), .B1(n4402), .B2(rd_idexe[1]), 
        .ZN(n7305) );
  AOI221_X1 U7679 ( .B1(n4083), .B2(rd_idexe[0]), .C1(n4402), .C2(rd_idexe[1]), 
        .A(n7305), .ZN(n7307) );
  XNOR2_X1 U7680 ( .A(rd_idexe[4]), .B(rs_id[4]), .ZN(n7306) );
  NAND4_X1 U7681 ( .A1(\ctrl_u/curr_exe[15] ), .A2(n7308), .A3(n7307), .A4(
        n7306), .ZN(n7310) );
  XOR2_X1 U7682 ( .A(n4370), .B(n4008), .Z(n7309) );
  AOI22_X1 U7683 ( .A1(\ctrl_u/curr_exe[0] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[0] ), .B2(n7337), .ZN(n7313) );
  INV_X1 U7684 ( .A(n7313), .ZN(\ctrl_u/next_exe[0] ) );
  AOI22_X1 U7685 ( .A1(\ctrl_u/curr_exe[10] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[10] ), .B2(n7337), .ZN(n7314) );
  INV_X1 U7686 ( .A(n7314), .ZN(\ctrl_u/next_exe[10] ) );
  AOI22_X1 U7687 ( .A1(\ctrl_u/curr_exe[11] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[11] ), .B2(n7337), .ZN(n7315) );
  INV_X1 U7688 ( .A(n7315), .ZN(\ctrl_u/next_exe[11] ) );
  AOI22_X1 U7689 ( .A1(\ctrl_u/curr_exe[12] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[12] ), .B2(n7337), .ZN(n7316) );
  INV_X1 U7690 ( .A(n7316), .ZN(\ctrl_u/next_exe[12] ) );
  AOI22_X1 U7691 ( .A1(\ctrl_u/curr_exe[13] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[13] ), .B2(n7337), .ZN(n7317) );
  INV_X1 U7692 ( .A(n7317), .ZN(\ctrl_u/next_exe[13] ) );
  AOI22_X1 U7693 ( .A1(\ctrl_u/curr_exe[14] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[14] ), .B2(n7337), .ZN(n7318) );
  INV_X1 U7694 ( .A(n7318), .ZN(\ctrl_u/next_exe[14] ) );
  AOI22_X1 U7695 ( .A1(\ctrl_u/curr_exe[16] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[16] ), .B2(n7337), .ZN(n7319) );
  INV_X1 U7696 ( .A(n7319), .ZN(\ctrl_u/next_exe[16] ) );
  AOI22_X1 U7697 ( .A1(\ctrl_u/curr_exe[19] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[19] ), .B2(n7337), .ZN(n7320) );
  INV_X1 U7698 ( .A(n7320), .ZN(\ctrl_u/next_exe[19] ) );
  AOI22_X1 U7699 ( .A1(\ctrl_u/curr_exe[1] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[1] ), .B2(n7337), .ZN(n7321) );
  INV_X1 U7700 ( .A(n7321), .ZN(\ctrl_u/next_exe[1] ) );
  AOI22_X1 U7701 ( .A1(\ctrl_u/curr_exe[20] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[20] ), .B2(n7337), .ZN(n7322) );
  INV_X1 U7702 ( .A(n7322), .ZN(\ctrl_u/next_exe[20] ) );
  AOI22_X1 U7703 ( .A1(alu_comp_sel[0]), .A2(n7338), .B1(\ctrl_u/curr_id[21] ), 
        .B2(n7337), .ZN(n7323) );
  INV_X1 U7704 ( .A(n7323), .ZN(\ctrl_u/next_exe[21] ) );
  AOI22_X1 U7705 ( .A1(op_sign_exe), .A2(n7338), .B1(\ctrl_u/curr_id[27] ), 
        .B2(n7337), .ZN(n7324) );
  INV_X1 U7706 ( .A(n7324), .ZN(\ctrl_u/next_exe[27] ) );
  AOI22_X1 U7707 ( .A1(op_type_exe[0]), .A2(n7338), .B1(\ctrl_u/curr_id[28] ), 
        .B2(n7337), .ZN(n7325) );
  INV_X1 U7708 ( .A(n7325), .ZN(\ctrl_u/next_exe[28] ) );
  AOI22_X1 U7709 ( .A1(log_type_exe[1]), .A2(n7338), .B1(\ctrl_u/curr_id[31] ), 
        .B2(n7337), .ZN(n7326) );
  INV_X1 U7710 ( .A(n7326), .ZN(\ctrl_u/next_exe[31] ) );
  AOI22_X1 U7711 ( .A1(log_type_exe[2]), .A2(n7338), .B1(\ctrl_u/curr_id[32] ), 
        .B2(n7337), .ZN(n7327) );
  INV_X1 U7712 ( .A(n7327), .ZN(\ctrl_u/next_exe[32] ) );
  AOI22_X1 U7713 ( .A1(log_type_exe[3]), .A2(n7338), .B1(\ctrl_u/curr_id[33] ), 
        .B2(n7337), .ZN(n7328) );
  INV_X1 U7714 ( .A(n7328), .ZN(\ctrl_u/next_exe[33] ) );
  AOI22_X1 U7715 ( .A1(shift_type_exe[2]), .A2(n7338), .B1(
        \ctrl_u/curr_id[36] ), .B2(n7337), .ZN(n7329) );
  INV_X1 U7716 ( .A(n7329), .ZN(\ctrl_u/next_exe[36] ) );
  AOI22_X1 U7717 ( .A1(sub_add_exe), .A2(n7338), .B1(\ctrl_u/curr_id[38] ), 
        .B2(n7337), .ZN(n7330) );
  INV_X1 U7718 ( .A(n7330), .ZN(\ctrl_u/next_exe[38] ) );
  AOI22_X1 U7719 ( .A1(\ctrl_u/curr_exe_39 ), .A2(n7338), .B1(
        \ctrl_u/curr_id[39] ), .B2(n7337), .ZN(n7331) );
  INV_X1 U7720 ( .A(n7331), .ZN(\ctrl_u/next_exe[39] ) );
  AOI22_X1 U7721 ( .A1(\ctrl_u/curr_exe_40 ), .A2(n7338), .B1(
        \ctrl_u/curr_id[40] ), .B2(n7337), .ZN(n7332) );
  INV_X1 U7722 ( .A(n7332), .ZN(\ctrl_u/next_exe[40] ) );
  AOI22_X1 U7723 ( .A1(\ctrl_u/curr_exe_41 ), .A2(n7338), .B1(
        \ctrl_u/curr_id[41] ), .B2(n7337), .ZN(n7333) );
  INV_X1 U7724 ( .A(n7333), .ZN(\ctrl_u/next_exe[41] ) );
  AOI22_X1 U7725 ( .A1(\ctrl_u/curr_exe[5] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[5] ), .B2(n7337), .ZN(n7334) );
  INV_X1 U7726 ( .A(n7334), .ZN(\ctrl_u/next_exe[5] ) );
  AOI22_X1 U7727 ( .A1(\ctrl_u/curr_exe[7] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[7] ), .B2(n7337), .ZN(n7335) );
  INV_X1 U7728 ( .A(n7335), .ZN(\ctrl_u/next_exe[7] ) );
  AOI22_X1 U7729 ( .A1(\ctrl_u/curr_exe[8] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[8] ), .B2(n7337), .ZN(n7336) );
  INV_X1 U7730 ( .A(n7336), .ZN(\ctrl_u/next_exe[8] ) );
  AOI22_X1 U7731 ( .A1(\ctrl_u/curr_exe[9] ), .A2(n7338), .B1(
        \ctrl_u/curr_id[9] ), .B2(n7337), .ZN(n7339) );
  INV_X1 U7732 ( .A(n7339), .ZN(\ctrl_u/next_exe[9] ) );
  NAND2_X1 U7733 ( .A1(n4209), .A2(n7370), .ZN(n7371) );
  NOR2_X1 U7734 ( .A1(n7371), .A2(\dp/npc_id_exe_int[6] ), .ZN(n7373) );
  NAND2_X1 U7735 ( .A1(n4210), .A2(n7373), .ZN(n7374) );
  NOR2_X1 U7736 ( .A1(n7374), .A2(\dp/npc_id_exe_int[8] ), .ZN(n7376) );
  NAND2_X1 U7737 ( .A1(n4217), .A2(n7376), .ZN(n7377) );
  NOR2_X1 U7738 ( .A1(n7377), .A2(\dp/npc_id_exe_int[10] ), .ZN(n7380) );
  NAND2_X1 U7739 ( .A1(n4218), .A2(n7380), .ZN(n7379) );
  NOR2_X1 U7740 ( .A1(n7379), .A2(\dp/npc_id_exe_int[12] ), .ZN(n7342) );
  AOI21_X1 U7741 ( .B1(n7379), .B2(\dp/npc_id_exe_int[12] ), .A(n7342), .ZN(
        n7341) );
  INV_X1 U7742 ( .A(n7341), .ZN(btb_cache_rw_address[10]) );
  NAND2_X1 U7743 ( .A1(n4226), .A2(n7342), .ZN(n7343) );
  OAI21_X1 U7744 ( .B1(n7342), .B2(n4226), .A(n7343), .ZN(
        btb_cache_rw_address[11]) );
  NOR2_X1 U7745 ( .A1(n7343), .A2(\dp/npc_id_exe_int[14] ), .ZN(n7345) );
  AOI21_X1 U7746 ( .B1(n7343), .B2(\dp/npc_id_exe_int[14] ), .A(n7345), .ZN(
        n7344) );
  INV_X1 U7747 ( .A(n7344), .ZN(btb_cache_rw_address[12]) );
  NAND2_X1 U7748 ( .A1(n4207), .A2(n7345), .ZN(n7346) );
  OAI21_X1 U7749 ( .B1(n7345), .B2(n4207), .A(n7346), .ZN(
        btb_cache_rw_address[13]) );
  NOR2_X1 U7750 ( .A1(n7346), .A2(\dp/npc_id_exe_int[16] ), .ZN(n7348) );
  AOI21_X1 U7751 ( .B1(n7346), .B2(\dp/npc_id_exe_int[16] ), .A(n7348), .ZN(
        n7347) );
  INV_X1 U7752 ( .A(n7347), .ZN(btb_cache_rw_address[14]) );
  NAND2_X1 U7753 ( .A1(\intadd_2/B[14] ), .A2(n7348), .ZN(n7349) );
  OAI21_X1 U7754 ( .B1(n7348), .B2(\intadd_2/B[14] ), .A(n7349), .ZN(
        btb_cache_rw_address[15]) );
  NOR2_X1 U7755 ( .A1(n7349), .A2(\dp/npc_id_exe_int[18] ), .ZN(n7351) );
  AOI21_X1 U7756 ( .B1(n7349), .B2(\dp/npc_id_exe_int[18] ), .A(n7351), .ZN(
        n7350) );
  INV_X1 U7757 ( .A(n7350), .ZN(btb_cache_rw_address[16]) );
  NAND2_X1 U7758 ( .A1(n4110), .A2(n7351), .ZN(n7352) );
  OAI21_X1 U7759 ( .B1(n7351), .B2(n4110), .A(n7352), .ZN(
        btb_cache_rw_address[17]) );
  NOR2_X1 U7760 ( .A1(n7352), .A2(\dp/npc_id_exe_int[20] ), .ZN(n7354) );
  AOI21_X1 U7761 ( .B1(n7352), .B2(\dp/npc_id_exe_int[20] ), .A(n7354), .ZN(
        n7353) );
  INV_X1 U7762 ( .A(n7353), .ZN(btb_cache_rw_address[18]) );
  NAND2_X1 U7763 ( .A1(n4101), .A2(n7354), .ZN(n7355) );
  OAI21_X1 U7764 ( .B1(n7354), .B2(n4101), .A(n7355), .ZN(
        btb_cache_rw_address[19]) );
  NOR2_X1 U7765 ( .A1(n7355), .A2(\dp/npc_id_exe_int[22] ), .ZN(n7357) );
  AOI21_X1 U7766 ( .B1(n7355), .B2(\dp/npc_id_exe_int[22] ), .A(n7357), .ZN(
        n7356) );
  INV_X1 U7767 ( .A(n7356), .ZN(btb_cache_rw_address[20]) );
  NAND2_X1 U7768 ( .A1(\intadd_2/B[20] ), .A2(n7357), .ZN(n7358) );
  OAI21_X1 U7769 ( .B1(n7357), .B2(\intadd_2/B[20] ), .A(n7358), .ZN(
        btb_cache_rw_address[21]) );
  NOR2_X1 U7770 ( .A1(n7358), .A2(\dp/npc_id_exe_int[24] ), .ZN(n7360) );
  AOI21_X1 U7771 ( .B1(n7358), .B2(\dp/npc_id_exe_int[24] ), .A(n7360), .ZN(
        n7359) );
  INV_X1 U7772 ( .A(n7359), .ZN(btb_cache_rw_address[22]) );
  NAND2_X1 U7773 ( .A1(n4137), .A2(n7360), .ZN(n7361) );
  OAI21_X1 U7774 ( .B1(n7360), .B2(n4137), .A(n7361), .ZN(
        btb_cache_rw_address[23]) );
  NOR2_X1 U7775 ( .A1(n7361), .A2(\dp/npc_id_exe_int[26] ), .ZN(n7363) );
  AOI21_X1 U7776 ( .B1(n7361), .B2(\dp/npc_id_exe_int[26] ), .A(n7363), .ZN(
        n7362) );
  INV_X1 U7777 ( .A(n7362), .ZN(btb_cache_rw_address[24]) );
  NAND2_X1 U7778 ( .A1(n4520), .A2(n7363), .ZN(n7364) );
  OAI21_X1 U7779 ( .B1(n7363), .B2(n4520), .A(n7364), .ZN(
        btb_cache_rw_address[25]) );
  NOR2_X1 U7780 ( .A1(n7364), .A2(\dp/npc_id_exe_int[28] ), .ZN(n7366) );
  AOI21_X1 U7781 ( .B1(n7364), .B2(\dp/npc_id_exe_int[28] ), .A(n7366), .ZN(
        n7365) );
  INV_X1 U7782 ( .A(n7365), .ZN(btb_cache_rw_address[26]) );
  NAND2_X1 U7783 ( .A1(n4536), .A2(n7366), .ZN(n7367) );
  OAI21_X1 U7784 ( .B1(n7366), .B2(n4536), .A(n7367), .ZN(
        btb_cache_rw_address[27]) );
  INV_X1 U7785 ( .A(n7367), .ZN(n7368) );
  NAND2_X1 U7786 ( .A1(n7368), .A2(n4519), .ZN(n7369) );
  OAI21_X1 U7787 ( .B1(n7368), .B2(n4519), .A(n7369), .ZN(
        btb_cache_rw_address[28]) );
  XNOR2_X1 U7788 ( .A(\dp/npc_id_exe_int[31] ), .B(n7369), .ZN(
        btb_cache_rw_address[29]) );
  OAI21_X1 U7789 ( .B1(n7370), .B2(n4209), .A(n7371), .ZN(
        btb_cache_rw_address[3]) );
  AOI21_X1 U7790 ( .B1(n7371), .B2(\dp/npc_id_exe_int[6] ), .A(n7373), .ZN(
        n7372) );
  INV_X1 U7791 ( .A(n7372), .ZN(btb_cache_rw_address[4]) );
  OAI21_X1 U7792 ( .B1(n7373), .B2(n4210), .A(n7374), .ZN(
        btb_cache_rw_address[5]) );
  AOI21_X1 U7793 ( .B1(n7374), .B2(\dp/npc_id_exe_int[8] ), .A(n7376), .ZN(
        n7375) );
  INV_X1 U7794 ( .A(n7375), .ZN(btb_cache_rw_address[6]) );
  OAI21_X1 U7795 ( .B1(n7376), .B2(n4217), .A(n7377), .ZN(
        btb_cache_rw_address[7]) );
  AOI21_X1 U7796 ( .B1(n7377), .B2(\dp/npc_id_exe_int[10] ), .A(n7380), .ZN(
        n7378) );
  INV_X1 U7797 ( .A(n7378), .ZN(btb_cache_rw_address[8]) );
  OAI21_X1 U7798 ( .B1(n7380), .B2(n4218), .A(n7379), .ZN(
        btb_cache_rw_address[9]) );
  NOR2_X1 U7800 ( .A1(n7428), .A2(n5229), .ZN(n7429) );
  AOI22_X1 U7801 ( .A1(n4021), .A2(n7429), .B1(n7428), .B2(rd[4]), .ZN(n1688)
         );
  NAND2_X1 U7802 ( .A1(rst_mem_wb_regs), .A2(en_cache_mem), .ZN(n7381) );
  AOI22_X1 U7803 ( .A1(\dp/cache_data_mem_wb_int[0] ), .A2(n7414), .B1(n7383), 
        .B2(\dp/cache_in_mem_int[0] ), .ZN(n1687) );
  AOI22_X1 U7804 ( .A1(\dp/cache_data_mem_wb_int[1] ), .A2(n7414), .B1(n7383), 
        .B2(\dp/cache_in_mem_int[1] ), .ZN(n1686) );
  AOI22_X1 U7805 ( .A1(\dp/cache_data_mem_wb_int[2] ), .A2(n7414), .B1(n7383), 
        .B2(\dp/cache_in_mem_int[2] ), .ZN(n1685) );
  AOI22_X1 U7806 ( .A1(\dp/cache_data_mem_wb_int[3] ), .A2(n7414), .B1(n7383), 
        .B2(\dp/cache_in_mem_int[3] ), .ZN(n1684) );
  AOI22_X1 U7807 ( .A1(\dp/cache_data_mem_wb_int[4] ), .A2(n7414), .B1(n7383), 
        .B2(\dp/cache_in_mem_int[4] ), .ZN(n1683) );
  AOI22_X1 U7808 ( .A1(\dp/cache_data_mem_wb_int[5] ), .A2(n7414), .B1(n7383), 
        .B2(\dp/cache_in_mem_int[5] ), .ZN(n1682) );
  AOI22_X1 U7809 ( .A1(\dp/cache_data_mem_wb_int[6] ), .A2(n7414), .B1(n7383), 
        .B2(\dp/cache_in_mem_int[6] ), .ZN(n1681) );
  AOI22_X1 U7810 ( .A1(\dp/cache_data_mem_wb_int[7] ), .A2(n7414), .B1(n7383), 
        .B2(\dp/cache_in_mem_int[7] ), .ZN(n1680) );
  NOR2_X1 U7811 ( .A1(ld_type_mem[0]), .A2(n4386), .ZN(n7382) );
  NAND4_X1 U7812 ( .A1(n7383), .A2(\dp/cache_in_mem_int[7] ), .A3(n7382), .A4(
        ld_sign_mem), .ZN(n7391) );
  AOI21_X1 U7813 ( .B1(n7396), .B2(dcache_data_in[8]), .A(n7394), .ZN(n7384)
         );
  AOI21_X1 U7814 ( .B1(n7396), .B2(dcache_data_in[9]), .A(n7394), .ZN(n7385)
         );
  AOI21_X1 U7815 ( .B1(n7396), .B2(dcache_data_in[10]), .A(n7394), .ZN(n7386)
         );
  AOI21_X1 U7816 ( .B1(n7396), .B2(dcache_data_in[11]), .A(n7394), .ZN(n7387)
         );
  AOI21_X1 U7817 ( .B1(n7396), .B2(dcache_data_in[12]), .A(n7394), .ZN(n7388)
         );
  AOI21_X1 U7818 ( .B1(n7396), .B2(dcache_data_in[13]), .A(n7394), .ZN(n7389)
         );
  AOI21_X1 U7819 ( .B1(n7396), .B2(dcache_data_in[14]), .A(n7394), .ZN(n7390)
         );
  NAND2_X1 U7820 ( .A1(n7396), .A2(dcache_data_in[15]), .ZN(n7393) );
  NAND2_X1 U7821 ( .A1(ld_type_mem[0]), .A2(n4386), .ZN(n7397) );
  NOR2_X1 U7822 ( .A1(n7393), .A2(n7397), .ZN(n7395) );
  AOI22_X1 U7823 ( .A1(\dp/cache_data_mem_wb_int[16] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[16]), .ZN(n7398) );
  NAND2_X1 U7824 ( .A1(n7416), .A2(n7398), .ZN(n3130) );
  AOI22_X1 U7825 ( .A1(\dp/cache_data_mem_wb_int[17] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[17]), .ZN(n7399) );
  NAND2_X1 U7826 ( .A1(n7416), .A2(n7399), .ZN(n3129) );
  AOI22_X1 U7827 ( .A1(\dp/cache_data_mem_wb_int[18] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[18]), .ZN(n7400) );
  NAND2_X1 U7828 ( .A1(n7416), .A2(n7400), .ZN(n3128) );
  AOI22_X1 U7829 ( .A1(\dp/cache_data_mem_wb_int[19] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[19]), .ZN(n7401) );
  NAND2_X1 U7830 ( .A1(n7416), .A2(n7401), .ZN(n3127) );
  AOI22_X1 U7831 ( .A1(\dp/cache_data_mem_wb_int[20] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[20]), .ZN(n7402) );
  NAND2_X1 U7832 ( .A1(n7416), .A2(n7402), .ZN(n3126) );
  AOI22_X1 U7833 ( .A1(\dp/cache_data_mem_wb_int[21] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[21]), .ZN(n7403) );
  NAND2_X1 U7834 ( .A1(n7416), .A2(n7403), .ZN(n3125) );
  AOI22_X1 U7835 ( .A1(\dp/cache_data_mem_wb_int[22] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[22]), .ZN(n7404) );
  NAND2_X1 U7836 ( .A1(n7416), .A2(n7404), .ZN(n3124) );
  AOI22_X1 U7837 ( .A1(\dp/cache_data_mem_wb_int[23] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[23]), .ZN(n7405) );
  NAND2_X1 U7838 ( .A1(n7416), .A2(n7405), .ZN(n3123) );
  AOI22_X1 U7839 ( .A1(\dp/cache_data_mem_wb_int[24] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[24]), .ZN(n7406) );
  NAND2_X1 U7840 ( .A1(n7416), .A2(n7406), .ZN(n3122) );
  AOI22_X1 U7841 ( .A1(\dp/cache_data_mem_wb_int[25] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[25]), .ZN(n7407) );
  NAND2_X1 U7842 ( .A1(n7416), .A2(n7407), .ZN(n3121) );
  AOI22_X1 U7843 ( .A1(\dp/cache_data_mem_wb_int[26] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[26]), .ZN(n7408) );
  NAND2_X1 U7844 ( .A1(n7416), .A2(n7408), .ZN(n3120) );
  AOI22_X1 U7845 ( .A1(\dp/cache_data_mem_wb_int[27] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[27]), .ZN(n7409) );
  NAND2_X1 U7846 ( .A1(n7416), .A2(n7409), .ZN(n3119) );
  AOI22_X1 U7847 ( .A1(\dp/cache_data_mem_wb_int[28] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[28]), .ZN(n7410) );
  NAND2_X1 U7848 ( .A1(n7416), .A2(n7410), .ZN(n3118) );
  AOI22_X1 U7849 ( .A1(\dp/cache_data_mem_wb_int[29] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[29]), .ZN(n7411) );
  NAND2_X1 U7850 ( .A1(n7416), .A2(n7411), .ZN(n3117) );
  AOI22_X1 U7851 ( .A1(\dp/cache_data_mem_wb_int[30] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[30]), .ZN(n7412) );
  NAND2_X1 U7852 ( .A1(n7416), .A2(n7412), .ZN(n3116) );
  AOI22_X1 U7853 ( .A1(\dp/cache_data_mem_wb_int[31] ), .A2(n7414), .B1(n7413), 
        .B2(dcache_data_in[31]), .ZN(n7415) );
  NAND2_X1 U7854 ( .A1(n7416), .A2(n7415), .ZN(n3115) );
  INV_X1 U7855 ( .A(evicted_cache_address[0]), .ZN(n7417) );
  OAI22_X1 U7856 ( .A1(n288), .A2(n3963), .B1(n7425), .B2(n7417), .ZN(n3112)
         );
  INV_X1 U7857 ( .A(evicted_cache_address[1]), .ZN(n7418) );
  OAI22_X1 U7858 ( .A1(n289), .A2(n3963), .B1(n7425), .B2(n7418), .ZN(n3111)
         );
  INV_X1 U7859 ( .A(evicted_cache_address[2]), .ZN(n7419) );
  OAI22_X1 U7860 ( .A1(n290), .A2(n3963), .B1(n7425), .B2(n7419), .ZN(n3110)
         );
  INV_X1 U7861 ( .A(evicted_cache_address[3]), .ZN(n7420) );
  OAI22_X1 U7862 ( .A1(n291), .A2(n3963), .B1(n7425), .B2(n7420), .ZN(n3109)
         );
  INV_X1 U7863 ( .A(evicted_cache_address[4]), .ZN(n7421) );
  OAI22_X1 U7864 ( .A1(n292), .A2(n3963), .B1(n7425), .B2(n7421), .ZN(n3108)
         );
  INV_X1 U7865 ( .A(evicted_cache_address[5]), .ZN(n7422) );
  OAI22_X1 U7866 ( .A1(n293), .A2(n3963), .B1(n7425), .B2(n7422), .ZN(n3107)
         );
  INV_X1 U7867 ( .A(evicted_cache_address[6]), .ZN(n7423) );
  OAI22_X1 U7868 ( .A1(n294), .A2(n3963), .B1(n7425), .B2(n7423), .ZN(n3106)
         );
  INV_X1 U7869 ( .A(evicted_cache_address[7]), .ZN(n7424) );
  OAI22_X1 U7870 ( .A1(n295), .A2(n3963), .B1(n7425), .B2(n7424), .ZN(n3105)
         );
  OAI22_X1 U7871 ( .A1(n299), .A2(n3963), .B1(n7425), .B2(n7500), .ZN(n3104)
         );
  OAI22_X1 U7872 ( .A1(n300), .A2(n3963), .B1(n7425), .B2(n7511), .ZN(n3103)
         );
  OAI22_X1 U7873 ( .A1(n301), .A2(n3963), .B1(n7425), .B2(n7522), .ZN(n3102)
         );
  OAI22_X1 U7874 ( .A1(n302), .A2(n3963), .B1(n7425), .B2(n7525), .ZN(n3101)
         );
  OAI22_X1 U7875 ( .A1(n303), .A2(n3963), .B1(n7425), .B2(n7526), .ZN(n3100)
         );
  OAI22_X1 U7876 ( .A1(n304), .A2(n3963), .B1(n7425), .B2(n7527), .ZN(n3099)
         );
  OAI22_X1 U7877 ( .A1(n305), .A2(n3963), .B1(n7425), .B2(n7528), .ZN(n3098)
         );
  OAI22_X1 U7878 ( .A1(n306), .A2(n3963), .B1(n7425), .B2(n7529), .ZN(n3097)
         );
  OAI22_X1 U7879 ( .A1(n307), .A2(n3963), .B1(n7425), .B2(n7530), .ZN(n3096)
         );
  OAI22_X1 U7880 ( .A1(n308), .A2(n3963), .B1(n7425), .B2(n7531), .ZN(n3095)
         );
  OAI22_X1 U7881 ( .A1(n309), .A2(n3963), .B1(n7425), .B2(n7501), .ZN(n3094)
         );
  OAI22_X1 U7882 ( .A1(n310), .A2(n3963), .B1(n7425), .B2(n7502), .ZN(n3093)
         );
  OAI22_X1 U7883 ( .A1(n311), .A2(n3963), .B1(n7425), .B2(n7503), .ZN(n3092)
         );
  OAI22_X1 U7884 ( .A1(n312), .A2(n3963), .B1(n7425), .B2(n7504), .ZN(n3091)
         );
  OAI22_X1 U7885 ( .A1(n313), .A2(n3963), .B1(n7425), .B2(n7505), .ZN(n3090)
         );
  OAI22_X1 U7886 ( .A1(n314), .A2(n3963), .B1(n7425), .B2(n7506), .ZN(n3089)
         );
  OAI22_X1 U7887 ( .A1(n315), .A2(n3963), .B1(n7425), .B2(n7507), .ZN(n3088)
         );
  OAI22_X1 U7888 ( .A1(n316), .A2(n3963), .B1(n7425), .B2(n7508), .ZN(n3087)
         );
  OAI22_X1 U7889 ( .A1(n317), .A2(n3963), .B1(n7425), .B2(n7509), .ZN(n3086)
         );
  OAI22_X1 U7890 ( .A1(n318), .A2(n3963), .B1(n7425), .B2(n7510), .ZN(n3085)
         );
  OAI22_X1 U7891 ( .A1(n319), .A2(n3963), .B1(n7425), .B2(n7512), .ZN(n3084)
         );
  OAI22_X1 U7892 ( .A1(n320), .A2(n3963), .B1(n7425), .B2(n7513), .ZN(n3083)
         );
  OAI22_X1 U7893 ( .A1(n321), .A2(n3963), .B1(n7425), .B2(n7514), .ZN(n3082)
         );
  OAI22_X1 U7894 ( .A1(n322), .A2(n3963), .B1(n7425), .B2(n7515), .ZN(n3081)
         );
  OAI22_X1 U7895 ( .A1(n323), .A2(n3963), .B1(n7425), .B2(n7516), .ZN(n3080)
         );
  OAI22_X1 U7896 ( .A1(n324), .A2(n3963), .B1(n7425), .B2(n7517), .ZN(n3079)
         );
  OAI22_X1 U7897 ( .A1(n325), .A2(n3963), .B1(n7425), .B2(n7518), .ZN(n3078)
         );
  OAI22_X1 U7898 ( .A1(n326), .A2(n3963), .B1(n7425), .B2(n7519), .ZN(n3077)
         );
  OAI22_X1 U7899 ( .A1(n327), .A2(n3963), .B1(n7425), .B2(n7520), .ZN(n3076)
         );
  OAI22_X1 U7900 ( .A1(n328), .A2(n3963), .B1(n7425), .B2(n7521), .ZN(n3075)
         );
  OAI22_X1 U7901 ( .A1(n329), .A2(n3963), .B1(n7425), .B2(n7523), .ZN(n3074)
         );
  OAI22_X1 U7902 ( .A1(n330), .A2(n3963), .B1(n7425), .B2(n7524), .ZN(n3073)
         );
  NAND2_X1 U7903 ( .A1(rst_mem_wb_regs), .A2(rst_exe_mem_regs), .ZN(n7442) );
  NOR2_X1 U7904 ( .A1(n7426), .A2(n7442), .ZN(n7427) );
  AOI22_X1 U7905 ( .A1(rd_idexe[0]), .A2(n7427), .B1(n7426), .B2(n4019), .ZN(
        n1606) );
  AOI22_X1 U7906 ( .A1(rd_idexe[1]), .A2(n7427), .B1(n7426), .B2(n3970), .ZN(
        n1605) );
  AOI22_X1 U7907 ( .A1(rd_idexe[2]), .A2(n7427), .B1(n7426), .B2(n4008), .ZN(
        n1604) );
  AOI22_X1 U7908 ( .A1(rd_idexe[3]), .A2(n7427), .B1(n7426), .B2(n4010), .ZN(
        n1603) );
  AOI22_X1 U7909 ( .A1(rd_idexe[4]), .A2(n7427), .B1(n7426), .B2(n4021), .ZN(
        n1600) );
  AOI22_X1 U7910 ( .A1(n4019), .A2(n7429), .B1(n7428), .B2(rd[0]), .ZN(n1599)
         );
  AOI22_X1 U7911 ( .A1(n3970), .A2(n7429), .B1(n7428), .B2(rd[1]), .ZN(n1598)
         );
  AOI22_X1 U7912 ( .A1(n4008), .A2(n7429), .B1(n7428), .B2(rd[2]), .ZN(n1597)
         );
  AOI22_X1 U7913 ( .A1(n4010), .A2(n7429), .B1(n7428), .B2(rd[3]), .ZN(n1594)
         );
  OAI22_X1 U7914 ( .A1(n4169), .A2(n5226), .B1(n7498), .B2(n4548), .ZN(n2786)
         );
  OAI22_X1 U7915 ( .A1(n4188), .A2(n5226), .B1(n7498), .B2(n4549), .ZN(n2785)
         );
  OAI22_X1 U7916 ( .A1(n7430), .A2(n5226), .B1(n5227), .B2(n4550), .ZN(n2784)
         );
  OAI22_X1 U7917 ( .A1(n4170), .A2(n5226), .B1(n5227), .B2(n4551), .ZN(n2783)
         );
  OAI22_X1 U7918 ( .A1(n4171), .A2(n5226), .B1(n7498), .B2(n4552), .ZN(n2782)
         );
  OAI22_X1 U7919 ( .A1(n4172), .A2(n5226), .B1(n5227), .B2(n4553), .ZN(n2781)
         );
  OAI22_X1 U7920 ( .A1(n4183), .A2(n5226), .B1(n5227), .B2(n4554), .ZN(n2780)
         );
  OAI22_X1 U7921 ( .A1(n4189), .A2(n5226), .B1(n5227), .B2(n4555), .ZN(n2779)
         );
  OAI22_X1 U7922 ( .A1(n7431), .A2(n5226), .B1(n5227), .B2(n4556), .ZN(n2778)
         );
  OAI22_X1 U7923 ( .A1(n4190), .A2(n5226), .B1(n7498), .B2(n4557), .ZN(n2777)
         );
  OAI22_X1 U7924 ( .A1(n4184), .A2(n5226), .B1(n5227), .B2(n4558), .ZN(n2776)
         );
  OAI22_X1 U7925 ( .A1(n4185), .A2(n5226), .B1(n5227), .B2(n4559), .ZN(n2775)
         );
  OAI22_X1 U7926 ( .A1(n4173), .A2(n5226), .B1(n7498), .B2(n4560), .ZN(n2774)
         );
  OAI22_X1 U7927 ( .A1(n4174), .A2(n5226), .B1(n5227), .B2(n4561), .ZN(n2773)
         );
  OAI22_X1 U7928 ( .A1(n7432), .A2(n5226), .B1(n5227), .B2(n4562), .ZN(n2772)
         );
  OAI22_X1 U7929 ( .A1(n4191), .A2(n5226), .B1(n7498), .B2(n4563), .ZN(n2771)
         );
  OAI22_X1 U7930 ( .A1(n4192), .A2(n5226), .B1(n7498), .B2(n4564), .ZN(n2770)
         );
  OAI22_X1 U7931 ( .A1(n4193), .A2(n5226), .B1(n5227), .B2(n4565), .ZN(n2769)
         );
  OAI22_X1 U7932 ( .A1(n7433), .A2(n5226), .B1(n7498), .B2(n4566), .ZN(n2768)
         );
  OAI22_X1 U7933 ( .A1(n4194), .A2(n5226), .B1(n7498), .B2(n4567), .ZN(n2767)
         );
  OAI22_X1 U7934 ( .A1(n4175), .A2(n5226), .B1(n7498), .B2(n4568), .ZN(n2766)
         );
  OAI22_X1 U7935 ( .A1(n4176), .A2(n5226), .B1(n7498), .B2(n4569), .ZN(n2765)
         );
  OAI22_X1 U7936 ( .A1(n4195), .A2(n5226), .B1(n7498), .B2(n4570), .ZN(n2764)
         );
  OAI22_X1 U7937 ( .A1(n4186), .A2(n5226), .B1(n7498), .B2(n4571), .ZN(n2763)
         );
  OAI22_X1 U7938 ( .A1(n4187), .A2(n5226), .B1(n7498), .B2(n4572), .ZN(n2762)
         );
  OAI22_X1 U7939 ( .A1(n4177), .A2(n5226), .B1(n7498), .B2(n4573), .ZN(n2761)
         );
  OAI22_X1 U7940 ( .A1(n4178), .A2(n5226), .B1(n7498), .B2(n4574), .ZN(n2760)
         );
  OAI22_X1 U7941 ( .A1(n4204), .A2(n5226), .B1(n7498), .B2(n4575), .ZN(n2759)
         );
  OAI22_X1 U7942 ( .A1(n7434), .A2(n5226), .B1(n7498), .B2(n4576), .ZN(n2758)
         );
  OAI22_X1 U7943 ( .A1(n4179), .A2(n5226), .B1(n7498), .B2(n4577), .ZN(n2757)
         );
  OAI22_X1 U7944 ( .A1(n7435), .A2(n5226), .B1(n7498), .B2(n4578), .ZN(n2756)
         );
  OAI22_X1 U7945 ( .A1(n681), .A2(n5226), .B1(n4539), .B2(n5227), .ZN(n2755)
         );
  NOR2_X1 U7946 ( .A1(b_selector_id), .A2(sign_ext_sel_id), .ZN(n7436) );
  OAI22_X1 U7947 ( .A1(n7437), .A2(n7440), .B1(n4089), .B2(n3942), .ZN(n2637)
         );
  OAI22_X1 U7948 ( .A1(n7438), .A2(n7440), .B1(n4095), .B2(n3938), .ZN(n2636)
         );
  INV_X1 U7949 ( .A(n7442), .ZN(n7441) );
  NAND2_X1 U7950 ( .A1(n7441), .A2(en_b_exe), .ZN(n7444) );
  INV_X1 U7951 ( .A(op_b_fw_sel_exe[1]), .ZN(n7443) );
  NOR3_X1 U7952 ( .A1(op_b_fw_sel_exe[0]), .A2(n7444), .A3(n7443), .ZN(n7491)
         );
  NAND2_X1 U7953 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[0] ), .ZN(n7447) );
  NAND2_X1 U7954 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[1] ), .ZN(n7448) );
  NAND2_X1 U7955 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[2] ), .ZN(n7449) );
  NAND2_X1 U7956 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[3] ), .ZN(n7450) );
  NAND2_X1 U7957 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[4] ), .ZN(n7451) );
  NAND2_X1 U7958 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[5] ), .ZN(n7452) );
  NAND2_X1 U7959 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[6] ), .ZN(n7453) );
  NAND2_X1 U7960 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[7] ), .ZN(n7454) );
  NAND2_X1 U7961 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[8] ), .ZN(n7455) );
  NAND2_X1 U7962 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[9] ), .ZN(n7456) );
  NAND2_X1 U7963 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[10] ), .ZN(n7457) );
  NAND2_X1 U7964 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[11] ), .ZN(n7458) );
  NAND2_X1 U7965 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[12] ), .ZN(n7459) );
  NAND2_X1 U7966 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[13] ), .ZN(n7460) );
  NAND2_X1 U7967 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[14] ), .ZN(n7461) );
  NAND2_X1 U7968 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[15] ), .ZN(n7462) );
  NAND2_X1 U7969 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[16] ), .ZN(n7463) );
  NAND2_X1 U7970 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[17] ), .ZN(n7464) );
  OAI211_X1 U7971 ( .C1(n7495), .C2(n4095), .A(n7465), .B(n7464), .ZN(n2604)
         );
  NAND2_X1 U7972 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[18] ), .ZN(n7466) );
  OAI211_X1 U7973 ( .C1(n7495), .C2(n4085), .A(n7467), .B(n7466), .ZN(n2603)
         );
  NAND2_X1 U7974 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[19] ), .ZN(n7468) );
  OAI211_X1 U7975 ( .C1(n7495), .C2(n4075), .A(n7469), .B(n7468), .ZN(n2602)
         );
  NAND2_X1 U7976 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[20] ), .ZN(n7470) );
  OAI211_X1 U7977 ( .C1(n7495), .C2(n4076), .A(n7471), .B(n7470), .ZN(n2601)
         );
  NAND2_X1 U7978 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[21] ), .ZN(n7472) );
  OAI211_X1 U7979 ( .C1(n7495), .C2(n4086), .A(n7473), .B(n7472), .ZN(n2600)
         );
  NAND2_X1 U7980 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[22] ), .ZN(n7474) );
  OAI211_X1 U7981 ( .C1(n7495), .C2(n4077), .A(n7475), .B(n7474), .ZN(n2599)
         );
  NAND2_X1 U7982 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[23] ), .ZN(n7476) );
  OAI211_X1 U7983 ( .C1(n7495), .C2(n4078), .A(n7477), .B(n7476), .ZN(n2598)
         );
  NAND2_X1 U7984 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[24] ), .ZN(n7478) );
  OAI211_X1 U7985 ( .C1(n7495), .C2(n4084), .A(n7479), .B(n7478), .ZN(n2597)
         );
  NAND2_X1 U7986 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[25] ), .ZN(n7480) );
  OAI211_X1 U7987 ( .C1(n7495), .C2(n4062), .A(n7481), .B(n7480), .ZN(n2596)
         );
  NAND2_X1 U7988 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[26] ), .ZN(n7482) );
  OAI211_X1 U7989 ( .C1(n7495), .C2(n4065), .A(n7483), .B(n7482), .ZN(n2595)
         );
  NAND2_X1 U7990 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[27] ), .ZN(n7484) );
  OAI211_X1 U7991 ( .C1(n7495), .C2(n4064), .A(n7485), .B(n7484), .ZN(n2594)
         );
  NAND2_X1 U7992 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[28] ), .ZN(n7486) );
  OAI211_X1 U7993 ( .C1(n7495), .C2(n4067), .A(n7487), .B(n7486), .ZN(n2593)
         );
  NAND2_X1 U7994 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[29] ), .ZN(n7488) );
  OAI211_X1 U7995 ( .C1(n7495), .C2(n4068), .A(n7489), .B(n7488), .ZN(n2592)
         );
  NAND2_X1 U7996 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[30] ), .ZN(n7490) );
  NAND2_X1 U7997 ( .A1(n7493), .A2(\dp/op_b_id_ex_int[31] ), .ZN(n7494) );
  OAI222_X1 U7998 ( .A1(n7499), .A2(n4196), .B1(n7497), .B2(n4089), .C1(n4587), 
        .C2(n5227), .ZN(n2573) );
  OAI222_X1 U7999 ( .A1(n7499), .A2(n4197), .B1(n7497), .B2(n4095), .C1(n4588), 
        .C2(n5227), .ZN(n2572) );
  OAI222_X1 U8000 ( .A1(n7499), .A2(n4198), .B1(n7497), .B2(n4085), .C1(n4589), 
        .C2(n5227), .ZN(n2571) );
  OAI222_X1 U8001 ( .A1(n7499), .A2(n4199), .B1(n7497), .B2(n4075), .C1(n4590), 
        .C2(n5227), .ZN(n2570) );
  OAI222_X1 U8002 ( .A1(n7499), .A2(n4200), .B1(n7497), .B2(n4076), .C1(n4591), 
        .C2(n5227), .ZN(n2569) );
  OAI222_X1 U8003 ( .A1(n7499), .A2(n4201), .B1(n7497), .B2(n4086), .C1(n4592), 
        .C2(n5227), .ZN(n2568) );
  OAI222_X1 U8004 ( .A1(n7499), .A2(n4202), .B1(n7497), .B2(n4077), .C1(n4593), 
        .C2(n5227), .ZN(n2567) );
  OAI222_X1 U8005 ( .A1(n7499), .A2(n4203), .B1(n7497), .B2(n4078), .C1(n4594), 
        .C2(n5227), .ZN(n2566) );
  OAI222_X1 U8006 ( .A1(n7499), .A2(n4530), .B1(n7497), .B2(n4084), .C1(n4112), 
        .C2(n5227), .ZN(n2565) );
  OAI222_X1 U8007 ( .A1(n7499), .A2(n4531), .B1(n7497), .B2(n4062), .C1(n4090), 
        .C2(n5227), .ZN(n2564) );
  OAI222_X1 U8008 ( .A1(n7499), .A2(n4532), .B1(n7497), .B2(n4065), .C1(n4091), 
        .C2(n5227), .ZN(n2563) );
  OAI222_X1 U8009 ( .A1(n7499), .A2(n4533), .B1(n7497), .B2(n4064), .C1(n4092), 
        .C2(n5227), .ZN(n2562) );
  OAI222_X1 U8010 ( .A1(n7499), .A2(n4534), .B1(n7497), .B2(n4067), .C1(n4093), 
        .C2(n5227), .ZN(n2561) );
  OAI222_X1 U8011 ( .A1(n7499), .A2(n4535), .B1(n7497), .B2(n4068), .C1(n4094), 
        .C2(n5227), .ZN(n2560) );
endmodule

