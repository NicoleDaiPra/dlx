library ieee;
use ieee.std_logic_1164.all;





-- ADD BITS TO ENABLE THE SAMPLING OF RS AND RT IN THE ID/EXE STAGE REGISTERS
-- BECAUSE OTHERWISE THE STALL UNIT USES THE WRONG REGISTERS (THE ONES OF ID) TO DETECT FORWARDING







package control_words is
	subtype cw_t is std_logic_vector(62 downto 0);
								   --  ID	       ID/EXE      EXE               E/M    MEM     M/W WB
	constant rtype_cw 		: cw_t := "000000000000000000000100000000000000001100011001000000000001000"; -- because the signals are determined using the func field
	constant bgez_bltz_cw 	: cw_t := "100000111101000000110011000000000010001101000000000000000000000";
	constant j_cw 			: cw_t := "010000101100000000110000000000000011101101000000000000000000000";
	constant jal_cw 		: cw_t := "010011100101000001110000000000000011101101011001000000001011100";
	constant beq_cw 		: cw_t := "100000111101000000110101000000000011001101000000000000000000000";
	constant bne_cw 		: cw_t := "100000111101000000110101000000000011011101000000000000000000000";
	constant blez_cw 		: cw_t := "100000111101000000110011000000000010001101000000000000000000000";
	constant bgtz_cw 		: cw_t := "100000111101000000110011000000000010111101000000000000000000000";
	constant addi_cw 		: cw_t := "100000111001000001000010000000000011111100011001000000001011100";
	constant addui_cw 		: cw_t := "100000011001000001000010000000000001111100011001000000001011100";
	constant subi_cw 		: cw_t := "100000111001000001000011000000000011111100011001000000001011100";
	constant subui_cw 		: cw_t := "100000011001000001000011000000000001111100011001000000001011100";
	constant andi_cw 		: cw_t := "100000011001000001000010000010001101111100011001000000001011100";
	constant ori_cw 		: cw_t := "100000011001000001000010000011101101111100011001000000001011100";
	constant xori_cw 		: cw_t := "100000011001000001000010000001101101111100011001000000001011100";
	constant beqz_cw 		: cw_t := "100000111101000000110011000000000011001101000000000000000000000";
	constant bnez_cw 		: cw_t := "100000111101000000110011000000000011011101000000000000000000000";
	constant slli_cw 		: cw_t := "100000011000010001000010001100001001111100011001000000001011100";
	constant srli_cw 		: cw_t := "100000011000010001000010001000001001111100011001000000001011100";
	constant srai_cw 		: cw_t := "100000011000010001000010010000001001111100011001000000001011100";
	constant seqi_cw 		: cw_t := "100000111001000001000011000000000011001000011001000000001011100";
	constant snei_cw 		: cw_t := "100000111001000001000011000000000011011010011001000000001011100";
	constant slti_cw 		: cw_t := "100000111001000001000011000000000010010010011001000000001011100";
	constant sgti_cw 		: cw_t := "100000111001000001000011000000000010110110011001000000001011100";
	constant slei_cw 		: cw_t := "100000111001000001000011000000000010000000011001000000001011100";
	constant sgei_cw 		: cw_t := "100000111001000001000011000000000010100100011001000000001011100";
	constant lb_cw			: cw_t := "100000111001000001000010000000000011111100011001100011000111110";
	constant lh_cw	 		: cw_t := "100000111001000001000010000000000011111100011001100010100111110";
	constant lw_cw	 		: cw_t := "100000111001000001000010000000000011111100011001100010000111110";
	constant lbu_cw 		: cw_t := "100000111001000001000010000000000011111100011001100001000111110";
	constant lhu_cw 		: cw_t := "100000111001000001000010000000000011111100011001100000100111110";
	constant sb_cw 			: cw_t := "100000111001000000001100000000000011111100011010011100010000000";
	constant sh_cw 			: cw_t := "100000111001000000001100000000000011111100011010011000010000000";
	constant sw_cw	 		: cw_t := "100000111001000000001100000000000011111100011010010100010000000";
	constant sltui_cw 		: cw_t := "100000111001000001000011000000000000010010011001000000001011100";
	constant sgtui_cw 		: cw_t := "100000111001000001000011000000000000110110011001000000001011100";
	constant sleui_cw 		: cw_t := "100000111001000001000011000000000000000000011001000000001011100";
	constant sgeui_cw 		: cw_t := "100000111001000001000011000000000000100100011001000000001011100";
end package control_words;