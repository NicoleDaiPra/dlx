library ieee;
use ieee.std_logic_1164.all;

package func_words is
	subtype fw_t is std_logic_vector(54 downto 0);
							   --  ID	        ID/EXE     EXE                E/M  MEM     M/W WB
	constant nop_func 	: fw_t	:= "00000001110 0010001000 000110000100000110 1100 0000000 101 100";
	constant sll_func 	: fw_t 	:= "00000001110 0010001000 000110000100000110 1100 0000000 101 100";
	constant srl_func 	: fw_t 	:= "00000001110 0010001000 000100000100000110 1100 0000000 101 100";
	constant sra_func 	: fw_t 	:= "00000001110 0010001000 001000000100000110 1100 0000000 101 100";
	constant jr_func 	: fw_t 	:= "01001101110 1000000000 000000000000000110 0000 0000000 000 000";
	constant jalr_func	: fw_t 	:= "01001101111 1000001001 000000000000000110 1101 0000001 101 100";
	constant mult_func 	: fw_t 	:= "00000001110 0100010000 000000000010000110 1000 0000000 100 001";
	constant mfhi_func 	: fw_t 	:= "00100001110 1000001000 000000000000000110 1100 0000000 101 100";
	constant mflo_func 	: fw_t 	:= "00010001110 1000001000 000000000000000110 1100 0000000 101 100";
	constant add_func 	: fw_t 	:= "00000001110 1000001000 000000000001000110 1100 0000000 101 100";
	constant addu_func 	: fw_t 	:= "00000001110 1000001000 000000000000000110 1100 0000000 101 100";
	constant sub_func 	: fw_t 	:= "00000001110 1000001000 100000000001000110 1100 0000000 101 100";
	constant subu_func 	: fw_t 	:= "00000001110 1000001000 100000000000000110 1100 0000000 101 100";
	constant and_func 	: fw_t 	:= "00000001110 1000001000 000001000110000110 1100 0000000 101 100";
	constant or_func 	: fw_t 	:= "00000001110 1000001000 000001110110000110 1100 0000000 101 100";
	constant xor_func 	: fw_t 	:= "00000001110 1000001000 000000110110000110 1100 0000000 101 100";
	constant seq_func 	: fw_t 	:= "00000001110 1000001000 100000000001000100 1100 0000000 101 100";
	constant sne_func 	: fw_t 	:= "00000001110 1000001000 100000000001000101 1100 0000000 101 100";
	constant slt_func 	: fw_t 	:= "00000001110 1000001000 100000000001000001 1100 0000000 101 100";
	constant sgt_func 	: fw_t 	:= "00000001110 1000001000 100000000001000011 1100 0000000 101 100";
	constant sle_func 	: fw_t 	:= "00000001110 1000001000 100000000001000000 1100 0000000 101 100";
	constant sge_func 	: fw_t 	:= "00000001110 1000001000 100000000001000010 1100 0000000 101 100";
	constant sltu_func 	: fw_t 	:= "00000001110 1000001000 100000000000000001 1100 0000000 101 100";
	constant sgtu_func 	: fw_t 	:= "00000001110 1000001000 100000000000000011 1100 0000000 101 100";
	constant sleu_func 	: fw_t 	:= "00000001110 1000001000 100000000000000000 1100 0000000 101 100";
	constant sgeu_func 	: fw_t 	:= "00000001110 1000001000 100000000000000010 1100 0000000 101 100";
end package func_words;